module lookuptable();
always@(negedge clk) begin
 case (w)
	12'b1_110_10000000 : r_w_inv <= 12'b1_111_01010101;
	12'b1_110_10000001 : r_w_inv <= 12'b1_111_01010101;
	12'b1_110_10000010 : r_w_inv <= 12'b1_111_01010101;
	12'b1_110_10000011 : r_w_inv <= 12'b1_111_01010100;
	12'b1_110_10000100 : r_w_inv <= 12'b1_111_01010100;
	12'b1_110_10000101 : r_w_inv <= 12'b1_111_01010011;
	12'b1_110_10000110 : r_w_inv <= 12'b1_111_01010011;
	12'b1_110_10000111 : r_w_inv <= 12'b1_111_01010010;
	12'b1_110_10001000 : r_w_inv <= 12'b1_111_01010010;
	12'b1_110_10001001 : r_w_inv <= 12'b1_111_01010001;
	12'b1_110_10001010 : r_w_inv <= 12'b1_111_01010001;
	12'b1_110_10001011 : r_w_inv <= 12'b1_111_01010000;
	12'b1_110_10001100 : r_w_inv <= 12'b1_111_01010000;
	12'b1_110_10001101 : r_w_inv <= 12'b1_111_01010000;
	12'b1_110_10001110 : r_w_inv <= 12'b1_111_01001111;
	12'b1_110_10001111 : r_w_inv <= 12'b1_111_01001111;
	12'b1_110_10010000 : r_w_inv <= 12'b1_111_01001110;
	12'b1_110_10010001 : r_w_inv <= 12'b1_111_01001110;
	12'b1_110_10010010 : r_w_inv <= 12'b1_111_01001101;
	12'b1_110_10010011 : r_w_inv <= 12'b1_111_01001101;
	12'b1_110_10010100 : r_w_inv <= 12'b1_111_01001100;
	12'b1_110_10010101 : r_w_inv <= 12'b1_111_01001100;
	12'b1_110_10010110 : r_w_inv <= 12'b1_111_01001011;
	12'b1_110_10010111 : r_w_inv <= 12'b1_111_01001011;
	12'b1_110_10011000 : r_w_inv <= 12'b1_111_01001010;
	12'b1_110_10011001 : r_w_inv <= 12'b1_111_01001010;
	12'b1_110_10011010 : r_w_inv <= 12'b1_111_01001001;
	12'b1_110_10011011 : r_w_inv <= 12'b1_111_01001001;
	12'b1_110_10011100 : r_w_inv <= 12'b1_111_01001000;
	12'b1_110_10011101 : r_w_inv <= 12'b1_111_01001000;
	12'b1_110_10011110 : r_w_inv <= 12'b1_111_01000111;
	12'b1_110_10011111 : r_w_inv <= 12'b1_111_01000110;
	12'b1_110_10100000 : r_w_inv <= 12'b1_111_01000110;
	12'b1_110_10100001 : r_w_inv <= 12'b1_111_01000110;
	12'b1_110_10100010 : r_w_inv <= 12'b1_111_01000101;
	12'b1_110_10100011 : r_w_inv <= 12'b1_111_01000100;
	12'b1_110_10100100 : r_w_inv <= 12'b1_111_01000100;
	12'b1_110_10100101 : r_w_inv <= 12'b1_111_01000011;
	12'b1_110_10100110 : r_w_inv <= 12'b1_111_01000011;
	12'b1_110_10100111 : r_w_inv <= 12'b1_111_01000010;
	12'b1_110_10101000 : r_w_inv <= 12'b1_111_01000010;
	12'b1_110_10101001 : r_w_inv <= 12'b1_111_01000001;
	12'b1_110_10101010 : r_w_inv <= 12'b1_111_01000001;
	12'b1_110_10101011 : r_w_inv <= 12'b1_111_01000000;
	12'b1_110_10101100 : r_w_inv <= 12'b1_111_01000000;
	12'b1_110_10101101 : r_w_inv <= 12'b1_111_00111111;
	12'b1_110_10101110 : r_w_inv <= 12'b1_111_00111110;
	12'b1_110_10101111 : r_w_inv <= 12'b1_111_00111110;
	12'b1_110_10110000 : r_w_inv <= 12'b1_111_00111101;
	12'b1_110_10110001 : r_w_inv <= 12'b1_111_00111101;
	12'b1_110_10110010 : r_w_inv <= 12'b1_111_00111100;
	12'b1_110_10110011 : r_w_inv <= 12'b1_111_00111011;
	12'b1_110_10110100 : r_w_inv <= 12'b1_111_00111011;
	12'b1_110_10110101 : r_w_inv <= 12'b1_111_00111010;
	12'b1_110_10110110 : r_w_inv <= 12'b1_111_00111010;
	12'b1_110_10110111 : r_w_inv <= 12'b1_111_00111001;
	12'b1_110_10111000 : r_w_inv <= 12'b1_111_00111000;
	12'b1_110_10111001 : r_w_inv <= 12'b1_111_00111000;
	12'b1_110_10111010 : r_w_inv <= 12'b1_111_00110111;
	12'b1_110_10111011 : r_w_inv <= 12'b1_111_00110111;
	12'b1_110_10111100 : r_w_inv <= 12'b1_111_00110110;
	12'b1_110_10111101 : r_w_inv <= 12'b1_111_00110101;
	12'b1_110_10111110 : r_w_inv <= 12'b1_111_00110101;
	12'b1_110_10111111 : r_w_inv <= 12'b1_111_00110100;
	12'b1_110_11000000 : r_w_inv <= 12'b1_111_00110011;
	12'b1_110_11000001 : r_w_inv <= 12'b1_111_00110011;
	12'b1_110_11000010 : r_w_inv <= 12'b1_111_00110010;
	12'b1_110_11000011 : r_w_inv <= 12'b1_111_00110010;
	12'b1_110_11000100 : r_w_inv <= 12'b1_111_00110001;
	12'b1_110_11000101 : r_w_inv <= 12'b1_111_00110000;
	12'b1_110_11000110 : r_w_inv <= 12'b1_111_00110000;
	12'b1_110_11000111 : r_w_inv <= 12'b1_111_00101111;
	12'b1_110_11001000 : r_w_inv <= 12'b1_111_00101110;
	12'b1_110_11001001 : r_w_inv <= 12'b1_111_00101101;
	12'b1_110_11001010 : r_w_inv <= 12'b1_111_00101101;
	12'b1_110_11001011 : r_w_inv <= 12'b1_111_00101100;
	12'b1_110_11001100 : r_w_inv <= 12'b1_111_00101100;
	12'b1_110_11001101 : r_w_inv <= 12'b1_111_00101011;
	12'b1_110_11001110 : r_w_inv <= 12'b1_111_00101010;
	12'b1_110_11001111 : r_w_inv <= 12'b1_111_00101001;
	12'b1_110_11010000 : r_w_inv <= 12'b1_111_00101001;
	12'b1_110_11010001 : r_w_inv <= 12'b1_111_00101000;
	12'b1_110_11010010 : r_w_inv <= 12'b1_111_00100111;
	12'b1_110_11010011 : r_w_inv <= 12'b1_111_00100110;
	12'b1_110_11010100 : r_w_inv <= 12'b1_111_00100110;
	12'b1_110_11010101 : r_w_inv <= 12'b1_111_00100101;
	12'b1_110_11010110 : r_w_inv <= 12'b1_111_00100100;
	12'b1_110_11010111 : r_w_inv <= 12'b1_111_00100100;
	12'b1_110_11011000 : r_w_inv <= 12'b1_111_00100011;
	12'b1_110_11011001 : r_w_inv <= 12'b1_111_00100010;
	12'b1_110_11011010 : r_w_inv <= 12'b1_111_00100001;
	12'b1_110_11011011 : r_w_inv <= 12'b1_111_00100001;
	12'b1_110_11011100 : r_w_inv <= 12'b1_111_00100000;
	12'b1_110_11011101 : r_w_inv <= 12'b1_111_00011111;
	12'b1_110_11011110 : r_w_inv <= 12'b1_111_00011110;
	12'b1_110_11011111 : r_w_inv <= 12'b1_111_00011101;
	12'b1_110_11100000 : r_w_inv <= 12'b1_111_00011101;
	12'b1_110_11100001 : r_w_inv <= 12'b1_111_00011100;
	12'b1_110_11100010 : r_w_inv <= 12'b1_111_00011011;
	12'b1_110_11100011 : r_w_inv <= 12'b1_111_00011010;
	12'b1_110_11100100 : r_w_inv <= 12'b1_111_00011010;
	12'b1_110_11100101 : r_w_inv <= 12'b1_111_00011001;
	12'b1_110_11100110 : r_w_inv <= 12'b1_111_00011000;
	12'b1_110_11100111 : r_w_inv <= 12'b1_111_00010111;
	12'b1_110_11101000 : r_w_inv <= 12'b1_111_00010110;
	12'b1_110_11101001 : r_w_inv <= 12'b1_111_00010101;
	12'b1_110_11101010 : r_w_inv <= 12'b1_111_00010100;
	12'b1_110_11101011 : r_w_inv <= 12'b1_111_00010100;
	12'b1_110_11101100 : r_w_inv <= 12'b1_111_00010011;
	12'b1_110_11101101 : r_w_inv <= 12'b1_111_00010010;
	12'b1_110_11101110 : r_w_inv <= 12'b1_111_00010001;
	12'b1_110_11101111 : r_w_inv <= 12'b1_111_00010000;
	12'b1_110_11110000 : r_w_inv <= 12'b1_111_00001111;
	12'b1_110_11110001 : r_w_inv <= 12'b1_111_00001110;
	12'b1_110_11110010 : r_w_inv <= 12'b1_111_00001110;
	12'b1_110_11110011 : r_w_inv <= 12'b1_111_00001101;
	12'b1_110_11110100 : r_w_inv <= 12'b1_111_00001100;
	12'b1_110_11110101 : r_w_inv <= 12'b1_111_00001011;
	12'b1_110_11110110 : r_w_inv <= 12'b1_111_00001010;
	12'b1_110_11110111 : r_w_inv <= 12'b1_111_00001001;
	12'b1_110_11111000 : r_w_inv <= 12'b1_111_00001000;
	12'b1_110_11111001 : r_w_inv <= 12'b1_111_00000111;
	12'b1_110_11111010 : r_w_inv <= 12'b1_111_00000110;
	12'b1_110_11111011 : r_w_inv <= 12'b1_111_00000101;
	12'b1_110_11111100 : r_w_inv <= 12'b1_111_00000100;
	12'b1_110_11111101 : r_w_inv <= 12'b1_111_00000011;
	12'b1_110_11111110 : r_w_inv <= 12'b1_111_00000010;
	12'b1_110_11111111 : r_w_inv <= 12'b1_111_00000001;
	12'b1_111_00000000 : r_w_inv <= 12'b1_111_00000000;
	12'b1_111_00000001 : r_w_inv <= 12'b1_110_11111111;
	12'b1_111_00000010 : r_w_inv <= 12'b1_110_11111110;
	12'b1_111_00000011 : r_w_inv <= 12'b1_110_11111101;
	12'b1_111_00000100 : r_w_inv <= 12'b1_110_11111100;
	12'b1_111_00000101 : r_w_inv <= 12'b1_110_11111011;
	12'b1_111_00000110 : r_w_inv <= 12'b1_110_11111010;
	12'b1_111_00000111 : r_w_inv <= 12'b1_110_11111001;
	12'b1_111_00001000 : r_w_inv <= 12'b1_110_11111000;
	12'b1_111_00001001 : r_w_inv <= 12'b1_110_11110111;
	12'b1_111_00001010 : r_w_inv <= 12'b1_110_11110110;
	12'b1_111_00001011 : r_w_inv <= 12'b1_110_11110101;
	12'b1_111_00001100 : r_w_inv <= 12'b1_110_11110100;
	12'b1_111_00001101 : r_w_inv <= 12'b1_110_11110011;
	12'b1_111_00001110 : r_w_inv <= 12'b1_110_11110010;
	12'b1_111_00001111 : r_w_inv <= 12'b1_110_11110001;
	12'b1_111_00010000 : r_w_inv <= 12'b1_110_11101111;
	12'b1_111_00010001 : r_w_inv <= 12'b1_110_11101110;
	12'b1_111_00010010 : r_w_inv <= 12'b1_110_11101101;
	12'b1_111_00010011 : r_w_inv <= 12'b1_110_11101100;
	12'b1_111_00010100 : r_w_inv <= 12'b1_110_11101011;
	12'b1_111_00010101 : r_w_inv <= 12'b1_110_11101001;
	12'b1_111_00010110 : r_w_inv <= 12'b1_110_11101001;
	12'b1_111_00010111 : r_w_inv <= 12'b1_110_11100111;
	12'b1_111_00011000 : r_w_inv <= 12'b1_110_11100110;
	12'b1_111_00011001 : r_w_inv <= 12'b1_110_11100101;
	12'b1_111_00011010 : r_w_inv <= 12'b1_110_11100100;
	12'b1_111_00011011 : r_w_inv <= 12'b1_110_11100010;
	12'b1_111_00011100 : r_w_inv <= 12'b1_110_11100001;
	12'b1_111_00011101 : r_w_inv <= 12'b1_110_11100000;
	12'b1_111_00011110 : r_w_inv <= 12'b1_110_11011110;
	12'b1_111_00011111 : r_w_inv <= 12'b1_110_11011101;
	12'b1_111_00100000 : r_w_inv <= 12'b1_110_11011100;
	12'b1_111_00100001 : r_w_inv <= 12'b1_110_11011011;
	12'b1_111_00100010 : r_w_inv <= 12'b1_110_11011001;
	12'b1_111_00100011 : r_w_inv <= 12'b1_110_11011000;
	12'b1_111_00100100 : r_w_inv <= 12'b1_110_11010111;
	12'b1_111_00100101 : r_w_inv <= 12'b1_110_11010101;
	12'b1_111_00100110 : r_w_inv <= 12'b1_110_11010100;
	12'b1_111_00100111 : r_w_inv <= 12'b1_110_11010010;
	12'b1_111_00101000 : r_w_inv <= 12'b1_110_11010001;
	12'b1_111_00101001 : r_w_inv <= 12'b1_110_11010000;
	12'b1_111_00101010 : r_w_inv <= 12'b1_110_11001110;
	12'b1_111_00101011 : r_w_inv <= 12'b1_110_11001101;
	12'b1_111_00101100 : r_w_inv <= 12'b1_110_11001100;
	12'b1_111_00101101 : r_w_inv <= 12'b1_110_11001010;
	12'b1_111_00101110 : r_w_inv <= 12'b1_110_11001001;
	12'b1_111_00101111 : r_w_inv <= 12'b1_110_11000111;
	12'b1_111_00110000 : r_w_inv <= 12'b1_110_11000110;
	12'b1_111_00110001 : r_w_inv <= 12'b1_110_11000100;
	12'b1_111_00110010 : r_w_inv <= 12'b1_110_11000010;
	12'b1_111_00110011 : r_w_inv <= 12'b1_110_11000001;
	12'b1_111_00110100 : r_w_inv <= 12'b1_110_10111111;
	12'b1_111_00110101 : r_w_inv <= 12'b1_110_10111110;
	12'b1_111_00110110 : r_w_inv <= 12'b1_110_10111100;
	12'b1_111_00110111 : r_w_inv <= 12'b1_110_10111011;
	12'b1_111_00111000 : r_w_inv <= 12'b1_110_10111001;
	12'b1_111_00111001 : r_w_inv <= 12'b1_110_10110111;
	12'b1_111_00111010 : r_w_inv <= 12'b1_110_10110110;
	12'b1_111_00111011 : r_w_inv <= 12'b1_110_10110100;
	12'b1_111_00111100 : r_w_inv <= 12'b1_110_10110010;
	12'b1_111_00111101 : r_w_inv <= 12'b1_110_10110000;
	12'b1_111_00111110 : r_w_inv <= 12'b1_110_10101111;
	12'b1_111_00111111 : r_w_inv <= 12'b1_110_10101101;
	12'b1_111_01000000 : r_w_inv <= 12'b1_110_10101011;
	12'b1_111_01000001 : r_w_inv <= 12'b1_110_10101010;
	12'b1_111_01000010 : r_w_inv <= 12'b1_110_10101000;
	12'b1_111_01000011 : r_w_inv <= 12'b1_110_10100110;
	12'b1_111_01000100 : r_w_inv <= 12'b1_110_10100100;
	12'b1_111_01000101 : r_w_inv <= 12'b1_110_10100010;
	12'b1_111_01000110 : r_w_inv <= 12'b1_110_10100000;
	12'b1_111_01000111 : r_w_inv <= 12'b1_110_10011110;
	12'b1_111_01001000 : r_w_inv <= 12'b1_110_10011100;
	12'b1_111_01001001 : r_w_inv <= 12'b1_110_10011010;
	12'b1_111_01001010 : r_w_inv <= 12'b1_110_10011000;
	12'b1_111_01001011 : r_w_inv <= 12'b1_110_10010110;
	12'b1_111_01001100 : r_w_inv <= 12'b1_110_10010101;
	12'b1_111_01001101 : r_w_inv <= 12'b1_110_10010011;
	12'b1_111_01001110 : r_w_inv <= 12'b1_110_10010001;
	12'b1_111_01001111 : r_w_inv <= 12'b1_110_10001111;
	12'b1_111_01010000 : r_w_inv <= 12'b1_110_10001100;
	12'b1_111_01010001 : r_w_inv <= 12'b1_110_10001010;
	12'b1_111_01010010 : r_w_inv <= 12'b1_110_10001000;
	12'b1_111_01010011 : r_w_inv <= 12'b1_110_10000110;
	12'b1_111_01010100 : r_w_inv <= 12'b1_110_10000100;
	12'b1_111_01010101 : r_w_inv <= 12'b1_110_10000001;
	12'b1_111_01010110 : r_w_inv <= 12'b1_110_10000000;
	12'b1_111_01010111 : r_w_inv <= 12'b1_110_01111101;
	12'b1_111_01011000 : r_w_inv <= 12'b1_110_01111011;
	12'b1_111_01011001 : r_w_inv <= 12'b1_110_01111001;
	12'b1_111_01011010 : r_w_inv <= 12'b1_110_01110110;
	12'b1_111_01011011 : r_w_inv <= 12'b1_110_01110100;
	12'b1_111_01011100 : r_w_inv <= 12'b1_110_01110001;
	12'b1_111_01011101 : r_w_inv <= 12'b1_110_01101111;
	12'b1_111_01011110 : r_w_inv <= 12'b1_110_01101100;
	12'b1_111_01011111 : r_w_inv <= 12'b1_110_01101010;
	12'b1_111_01100000 : r_w_inv <= 12'b1_110_01100111;
	12'b1_111_01100001 : r_w_inv <= 12'b1_110_01100101;
	12'b1_111_01100010 : r_w_inv <= 12'b1_110_01100010;
	12'b1_111_01100011 : r_w_inv <= 12'b1_110_01100000;
	12'b1_111_01100100 : r_w_inv <= 12'b1_110_01011101;
	12'b1_111_01100101 : r_w_inv <= 12'b1_110_01011010;
	12'b1_111_01100110 : r_w_inv <= 12'b1_110_01010111;
	12'b1_111_01100111 : r_w_inv <= 12'b1_110_01010101;
	12'b1_111_01101000 : r_w_inv <= 12'b1_110_01010010;
	12'b1_111_01101001 : r_w_inv <= 12'b1_110_01001111;
	12'b1_111_01101010 : r_w_inv <= 12'b1_110_01001100;
	12'b1_111_01101011 : r_w_inv <= 12'b1_110_01001001;
	12'b1_111_01101100 : r_w_inv <= 12'b1_110_01000111;
	12'b1_111_01101101 : r_w_inv <= 12'b1_110_01000100;
	12'b1_111_01101110 : r_w_inv <= 12'b1_110_01000000;
	12'b1_111_01101111 : r_w_inv <= 12'b1_110_00111101;
	12'b1_111_01110000 : r_w_inv <= 12'b1_110_00111010;
	12'b1_111_01110001 : r_w_inv <= 12'b1_110_00110111;
	12'b1_111_01110010 : r_w_inv <= 12'b1_110_00110100;
	12'b1_111_01110011 : r_w_inv <= 12'b1_110_00110000;
	12'b1_111_01110100 : r_w_inv <= 12'b1_110_00101101;
	12'b1_111_01110101 : r_w_inv <= 12'b1_110_00101001;
	12'b1_111_01110110 : r_w_inv <= 12'b1_110_00100111;
	12'b1_111_01110111 : r_w_inv <= 12'b1_110_00100011;
	12'b1_111_01111000 : r_w_inv <= 12'b1_110_00100000;
	12'b1_111_01111001 : r_w_inv <= 12'b1_110_00011100;
	12'b1_111_01111010 : r_w_inv <= 12'b1_110_00011000;
	12'b1_111_01111011 : r_w_inv <= 12'b1_110_00010101;
	12'b1_111_01111100 : r_w_inv <= 12'b1_110_00010001;
	12'b1_111_01111101 : r_w_inv <= 12'b1_110_00001101;
	12'b1_111_01111110 : r_w_inv <= 12'b1_110_00001001;
	12'b1_111_01111111 : r_w_inv <= 12'b1_110_00000101;
	12'b1_111_10000000 : r_w_inv <= 12'b1_110_00000001;
	12'b1_111_10000001 : r_w_inv <= 12'b1_101_11111110;
	12'b1_111_10000010 : r_w_inv <= 12'b1_101_11111010;
	12'b1_111_10000011 : r_w_inv <= 12'b1_101_11110110;
	12'b1_111_10000100 : r_w_inv <= 12'b1_101_11110001;
	12'b1_111_10000101 : r_w_inv <= 12'b1_101_11101101;
	12'b1_111_10000110 : r_w_inv <= 12'b1_101_11101000;
	12'b1_111_10000111 : r_w_inv <= 12'b1_101_11100100;
	12'b1_111_10001000 : r_w_inv <= 12'b1_101_11011111;
	12'b1_111_10001001 : r_w_inv <= 12'b1_101_11011011;
	12'b1_111_10001010 : r_w_inv <= 12'b1_101_11010110;
	12'b1_111_10001011 : r_w_inv <= 12'b1_101_11010001;
	12'b1_111_10001100 : r_w_inv <= 12'b1_101_11001101;
	12'b1_111_10001101 : r_w_inv <= 12'b1_101_11001000;
	12'b1_111_10001110 : r_w_inv <= 12'b1_101_11000011;
	12'b1_111_10001111 : r_w_inv <= 12'b1_101_10111110;
	12'b1_111_10010000 : r_w_inv <= 12'b1_101_10111001;
	12'b1_111_10010001 : r_w_inv <= 12'b1_101_10110011;
	12'b1_111_10010010 : r_w_inv <= 12'b1_101_10101110;
	12'b1_111_10010011 : r_w_inv <= 12'b1_101_10101000;
	12'b1_111_10010100 : r_w_inv <= 12'b1_101_10100011;
	12'b1_111_10010101 : r_w_inv <= 12'b1_101_10011101;
	12'b1_111_10010110 : r_w_inv <= 12'b1_101_10011001;
	12'b1_111_10010111 : r_w_inv <= 12'b1_101_10010011;
	12'b1_111_10011000 : r_w_inv <= 12'b1_101_10001101;
	12'b1_111_10011001 : r_w_inv <= 12'b1_101_10000110;
	12'b1_111_10011010 : r_w_inv <= 12'b1_101_10000000;
	12'b1_111_10011011 : r_w_inv <= 12'b1_101_01111010;
	12'b1_111_10011100 : r_w_inv <= 12'b1_101_01110011;
	12'b1_111_10011101 : r_w_inv <= 12'b1_101_01101100;
	12'b1_111_10011110 : r_w_inv <= 12'b1_101_01100101;
	12'b1_111_10011111 : r_w_inv <= 12'b1_101_01011110;
	12'b1_111_10100000 : r_w_inv <= 12'b1_101_01010111;
	12'b1_111_10100001 : r_w_inv <= 12'b1_101_01010010;
	12'b1_111_10100010 : r_w_inv <= 12'b1_101_01001010;
	12'b1_111_10100011 : r_w_inv <= 12'b1_101_01000011;
	12'b1_111_10100100 : r_w_inv <= 12'b1_101_00111011;
	12'b1_111_10100101 : r_w_inv <= 12'b1_101_00110011;
	12'b1_111_10100110 : r_w_inv <= 12'b1_101_00101011;
	12'b1_111_10100111 : r_w_inv <= 12'b1_101_00100010;
	12'b1_111_10101000 : r_w_inv <= 12'b1_101_00011010;
	12'b1_111_10101001 : r_w_inv <= 12'b1_101_00010001;
	12'b1_111_10101010 : r_w_inv <= 12'b1_101_00001000;
	12'b1_111_10101011 : r_w_inv <= 12'b1_100_11111111;
	12'b1_111_10101100 : r_w_inv <= 12'b1_100_11111000;
	12'b1_111_10101101 : r_w_inv <= 12'b1_100_11101111;
	12'b1_111_10101110 : r_w_inv <= 12'b1_100_11100101;
	12'b1_111_10101111 : r_w_inv <= 12'b1_100_11011011;
	12'b1_111_10110000 : r_w_inv <= 12'b1_100_11010001;
	12'b1_111_10110001 : r_w_inv <= 12'b1_100_11000110;
	12'b1_111_10110010 : r_w_inv <= 12'b1_100_10111011;
	12'b1_111_10110011 : r_w_inv <= 12'b1_100_10110000;
	12'b1_111_10110100 : r_w_inv <= 12'b1_100_10100101;
	12'b1_111_10110101 : r_w_inv <= 12'b1_100_10011001;
	12'b1_111_10110110 : r_w_inv <= 12'b1_100_10010000;
	12'b1_111_10110111 : r_w_inv <= 12'b1_100_10000100;
	12'b1_111_10111000 : r_w_inv <= 12'b1_100_01110111;
	12'b1_111_10111001 : r_w_inv <= 12'b1_100_01101010;
	12'b1_111_10111010 : r_w_inv <= 12'b1_100_01011101;
	12'b1_111_10111011 : r_w_inv <= 12'b1_100_01001111;
	12'b1_111_10111100 : r_w_inv <= 12'b1_100_01000001;
	12'b1_111_10111101 : r_w_inv <= 12'b1_100_00110011;
	12'b1_111_10111110 : r_w_inv <= 12'b1_100_00100100;
	12'b1_111_10111111 : r_w_inv <= 12'b1_100_00010100;
	12'b1_111_11000000 : r_w_inv <= 12'b1_100_00000100;
	12'b1_111_11000001 : r_w_inv <= 12'b1_011_11111000;
	12'b1_111_11000010 : r_w_inv <= 12'b1_011_11100111;
	12'b1_111_11000011 : r_w_inv <= 12'b1_011_11010101;
	12'b1_111_11000100 : r_w_inv <= 12'b1_011_11000011;
	12'b1_111_11000101 : r_w_inv <= 12'b1_011_10110001;
	12'b1_111_11000110 : r_w_inv <= 12'b1_011_10011101;
	12'b1_111_11000111 : r_w_inv <= 12'b1_011_10001001;
	12'b1_111_11001000 : r_w_inv <= 12'b1_011_01110100;
	12'b1_111_11001001 : r_w_inv <= 12'b1_011_01011111;
	12'b1_111_11001010 : r_w_inv <= 12'b1_011_01001000;
	12'b1_111_11001011 : r_w_inv <= 12'b1_011_00110001;
	12'b1_111_11001100 : r_w_inv <= 12'b1_011_00011111;
	12'b1_111_11001101 : r_w_inv <= 12'b1_011_00000110;
	12'b1_111_11001110 : r_w_inv <= 12'b1_010_11101101;
	12'b1_111_11001111 : r_w_inv <= 12'b1_010_11010010;
	12'b1_111_11010000 : r_w_inv <= 12'b1_010_10110110;
	12'b1_111_11010001 : r_w_inv <= 12'b1_010_10011000;
	12'b1_111_11010010 : r_w_inv <= 12'b1_010_01111010;
	12'b1_111_11010011 : r_w_inv <= 12'b1_010_01011010;
	12'b1_111_11010100 : r_w_inv <= 12'b1_010_00111000;
	12'b1_111_11010101 : r_w_inv <= 12'b1_010_00010101;
	12'b1_111_11010110 : r_w_inv <= 12'b1_001_11111010;
	12'b1_111_11010111 : r_w_inv <= 12'b1_001_11010100;
	12'b1_111_11011000 : r_w_inv <= 12'b1_001_10101100;
	12'b1_111_11011001 : r_w_inv <= 12'b1_001_10000010;
	12'b1_111_11011010 : r_w_inv <= 12'b1_001_01010101;
	12'b1_111_11011011 : r_w_inv <= 12'b1_001_00100111;
	12'b1_111_11011100 : r_w_inv <= 12'b1_000_11110101;
	12'b1_111_11011101 : r_w_inv <= 12'b1_000_11000001;
	12'b1_111_11011110 : r_w_inv <= 12'b1_000_10001010;
	12'b1_111_11011111 : r_w_inv <= 12'b1_000_01001111;
	12'b1_111_11100000 : r_w_inv <= 12'b1_000_00010000;
	12'b1_111_11100001 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11100010 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11100011 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11100100 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11100101 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11100110 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11100111 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11101000 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11101001 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11101010 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11101011 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11101100 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11101101 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11101110 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11101111 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11110000 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11110001 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11110010 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11110011 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11110100 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11110101 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11110110 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11110111 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11111000 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11111001 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11111010 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11111011 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11111100 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11111101 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11111110 : r_w_inv <= 12'b1_000_00000000;
	12'b1_111_11111111 : r_w_inv <= 12'b1_000_00000000;
	12'b0_000_00000000 : r_w_inv <= 12'b1_000_00000000;
	12'b0_000_00000001 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00000010 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00000011 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00000100 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00000101 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00000110 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00000111 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00001000 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00001001 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00001010 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00001011 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00001100 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00001101 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00001110 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00001111 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00010000 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00010001 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00010010 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00010011 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00010100 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00010101 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00010110 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00010111 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00011000 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00011001 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00011010 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00011011 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00011100 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00011101 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00011110 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00011111 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00100000 : r_w_inv <= 12'b0_111_11111111;
	12'b0_000_00100001 : r_w_inv <= 12'b0_111_11010000;
	12'b0_000_00100010 : r_w_inv <= 12'b0_111_10010011;
	12'b0_000_00100011 : r_w_inv <= 12'b0_111_01011010;
	12'b0_000_00100100 : r_w_inv <= 12'b0_111_00100101;
	12'b0_000_00100101 : r_w_inv <= 12'b0_110_11110010;
	12'b0_000_00100110 : r_w_inv <= 12'b0_110_11000010;
	12'b0_000_00100111 : r_w_inv <= 12'b0_110_10010100;
	12'b0_000_00101000 : r_w_inv <= 12'b0_110_01101001;
	12'b0_000_00101001 : r_w_inv <= 12'b0_110_01000000;
	12'b0_000_00101010 : r_w_inv <= 12'b0_110_00011001;
	12'b0_000_00101011 : r_w_inv <= 12'b0_101_11110100;
	12'b0_000_00101100 : r_w_inv <= 12'b0_101_11011001;
	12'b0_000_00101101 : r_w_inv <= 12'b0_101_10110111;
	12'b0_000_00101110 : r_w_inv <= 12'b0_101_10010110;
	12'b0_000_00101111 : r_w_inv <= 12'b0_101_01110111;
	12'b0_000_00110000 : r_w_inv <= 12'b0_101_01011001;
	12'b0_000_00110001 : r_w_inv <= 12'b0_101_00111100;
	12'b0_000_00110010 : r_w_inv <= 12'b0_101_00100001;
	12'b0_000_00110011 : r_w_inv <= 12'b0_101_00000110;
	12'b0_000_00110100 : r_w_inv <= 12'b0_100_11101101;
	12'b0_000_00110101 : r_w_inv <= 12'b0_100_11010101;
	12'b0_000_00110110 : r_w_inv <= 12'b0_100_11000011;
	12'b0_000_00110111 : r_w_inv <= 12'b0_100_10101100;
	12'b0_000_00111000 : r_w_inv <= 12'b0_100_10010110;
	12'b0_000_00111001 : r_w_inv <= 12'b0_100_10000001;
	12'b0_000_00111010 : r_w_inv <= 12'b0_100_01101101;
	12'b0_000_00111011 : r_w_inv <= 12'b0_100_01011001;
	12'b0_000_00111100 : r_w_inv <= 12'b0_100_01000110;
	12'b0_000_00111101 : r_w_inv <= 12'b0_100_00110100;
	12'b0_000_00111110 : r_w_inv <= 12'b0_100_00100010;
	12'b0_000_00111111 : r_w_inv <= 12'b0_100_00010001;
	12'b0_000_01000000 : r_w_inv <= 12'b0_100_00000000;
	12'b0_000_01000001 : r_w_inv <= 12'b0_011_11110100;
	12'b0_000_01000010 : r_w_inv <= 12'b0_011_11100100;
	12'b0_000_01000011 : r_w_inv <= 12'b0_011_11010101;
	12'b0_000_01000100 : r_w_inv <= 12'b0_011_11000110;
	12'b0_000_01000101 : r_w_inv <= 12'b0_011_10111000;
	12'b0_000_01000110 : r_w_inv <= 12'b0_011_10101010;
	12'b0_000_01000111 : r_w_inv <= 12'b0_011_10011100;
	12'b0_000_01001000 : r_w_inv <= 12'b0_011_10001111;
	12'b0_000_01001001 : r_w_inv <= 12'b0_011_10000010;
	12'b0_000_01001010 : r_w_inv <= 12'b0_011_01110110;
	12'b0_000_01001011 : r_w_inv <= 12'b0_011_01101010;
	12'b0_000_01001100 : r_w_inv <= 12'b0_011_01100001;
	12'b0_000_01001101 : r_w_inv <= 12'b0_011_01010101;
	12'b0_000_01001110 : r_w_inv <= 12'b0_011_01001010;
	12'b0_000_01001111 : r_w_inv <= 12'b0_011_00111111;
	12'b0_000_01010000 : r_w_inv <= 12'b0_011_00110101;
	12'b0_000_01010001 : r_w_inv <= 12'b0_011_00101010;
	12'b0_000_01010010 : r_w_inv <= 12'b0_011_00100000;
	12'b0_000_01010011 : r_w_inv <= 12'b0_011_00010110;
	12'b0_000_01010100 : r_w_inv <= 12'b0_011_00001100;
	12'b0_000_01010101 : r_w_inv <= 12'b0_011_00000011;
	12'b0_000_01010110 : r_w_inv <= 12'b0_010_11111100;
	12'b0_000_01010111 : r_w_inv <= 12'b0_010_11110011;
	12'b0_000_01011000 : r_w_inv <= 12'b0_010_11101010;
	12'b0_000_01011001 : r_w_inv <= 12'b0_010_11100010;
	12'b0_000_01011010 : r_w_inv <= 12'b0_010_11011001;
	12'b0_000_01011011 : r_w_inv <= 12'b0_010_11010001;
	12'b0_000_01011100 : r_w_inv <= 12'b0_010_11001001;
	12'b0_000_01011101 : r_w_inv <= 12'b0_010_11000001;
	12'b0_000_01011110 : r_w_inv <= 12'b0_010_10111010;
	12'b0_000_01011111 : r_w_inv <= 12'b0_010_10110010;
	12'b0_000_01100000 : r_w_inv <= 12'b0_010_10101011;
	12'b0_000_01100001 : r_w_inv <= 12'b0_010_10100101;
	12'b0_000_01100010 : r_w_inv <= 12'b0_010_10011110;
	12'b0_000_01100011 : r_w_inv <= 12'b0_010_10010111;
	12'b0_000_01100100 : r_w_inv <= 12'b0_010_10010000;
	12'b0_000_01100101 : r_w_inv <= 12'b0_010_10001010;
	12'b0_000_01100110 : r_w_inv <= 12'b0_010_10000011;
	12'b0_000_01100111 : r_w_inv <= 12'b0_010_01111101;
	12'b0_000_01101000 : r_w_inv <= 12'b0_010_01110111;
	12'b0_000_01101001 : r_w_inv <= 12'b0_010_01110000;
	12'b0_000_01101010 : r_w_inv <= 12'b0_010_01101010;
	12'b0_000_01101011 : r_w_inv <= 12'b0_010_01100100;
	12'b0_000_01101100 : r_w_inv <= 12'b0_010_01100000;
	12'b0_000_01101101 : r_w_inv <= 12'b0_010_01011010;
	12'b0_000_01101110 : r_w_inv <= 12'b0_010_01010101;
	12'b0_000_01101111 : r_w_inv <= 12'b0_010_01001111;
	12'b0_000_01110000 : r_w_inv <= 12'b0_010_01001010;
	12'b0_000_01110001 : r_w_inv <= 12'b0_010_01000100;
	12'b0_000_01110010 : r_w_inv <= 12'b0_010_00111111;
	12'b0_000_01110011 : r_w_inv <= 12'b0_010_00111010;
	12'b0_000_01110100 : r_w_inv <= 12'b0_010_00110101;
	12'b0_000_01110101 : r_w_inv <= 12'b0_010_00110000;
	12'b0_000_01110110 : r_w_inv <= 12'b0_010_00101101;
	12'b0_000_01110111 : r_w_inv <= 12'b0_010_00101000;
	12'b0_000_01111000 : r_w_inv <= 12'b0_010_00100011;
	12'b0_000_01111001 : r_w_inv <= 12'b0_010_00011110;
	12'b0_000_01111010 : r_w_inv <= 12'b0_010_00011010;
	12'b0_000_01111011 : r_w_inv <= 12'b0_010_00010101;
	12'b0_000_01111100 : r_w_inv <= 12'b0_010_00010001;
	12'b0_000_01111101 : r_w_inv <= 12'b0_010_00001101;
	12'b0_000_01111110 : r_w_inv <= 12'b0_010_00001000;
	12'b0_000_01111111 : r_w_inv <= 12'b0_010_00000100;
	12'b0_000_10000000 : r_w_inv <= 12'b0_010_00000000;
	12'b0_000_10000001 : r_w_inv <= 12'b0_001_11111101;
	12'b0_000_10000010 : r_w_inv <= 12'b0_001_11111001;
	12'b0_000_10000011 : r_w_inv <= 12'b0_001_11110101;
	12'b0_000_10000100 : r_w_inv <= 12'b0_001_11110001;
	12'b0_000_10000101 : r_w_inv <= 12'b0_001_11101101;
	12'b0_000_10000110 : r_w_inv <= 12'b0_001_11101001;
	12'b0_000_10000111 : r_w_inv <= 12'b0_001_11100110;
	12'b0_000_10001000 : r_w_inv <= 12'b0_001_11100010;
	12'b0_000_10001001 : r_w_inv <= 12'b0_001_11011111;
	12'b0_000_10001010 : r_w_inv <= 12'b0_001_11011011;
	12'b0_000_10001011 : r_w_inv <= 12'b0_001_11010111;
	12'b0_000_10001100 : r_w_inv <= 12'b0_001_11010101;
	12'b0_000_10001101 : r_w_inv <= 12'b0_001_11010001;
	12'b0_000_10001110 : r_w_inv <= 12'b0_001_11001110;
	12'b0_000_10001111 : r_w_inv <= 12'b0_001_11001011;
	12'b0_000_10010000 : r_w_inv <= 12'b0_001_11001000;
	12'b0_000_10010001 : r_w_inv <= 12'b0_001_11000100;
	12'b0_000_10010010 : r_w_inv <= 12'b0_001_11000001;
	12'b0_000_10010011 : r_w_inv <= 12'b0_001_10111110;
	12'b0_000_10010100 : r_w_inv <= 12'b0_001_10111011;
	12'b0_000_10010101 : r_w_inv <= 12'b0_001_10111000;
	12'b0_000_10010110 : r_w_inv <= 12'b0_001_10110110;
	12'b0_000_10010111 : r_w_inv <= 12'b0_001_10110011;
	12'b0_000_10011000 : r_w_inv <= 12'b0_001_10110000;
	12'b0_000_10011001 : r_w_inv <= 12'b0_001_10101101;
	12'b0_000_10011010 : r_w_inv <= 12'b0_001_10101010;
	12'b0_000_10011011 : r_w_inv <= 12'b0_001_10100111;
	12'b0_000_10011100 : r_w_inv <= 12'b0_001_10100100;
	12'b0_000_10011101 : r_w_inv <= 12'b0_001_10100010;
	12'b0_000_10011110 : r_w_inv <= 12'b0_001_10011111;
	12'b0_000_10011111 : r_w_inv <= 12'b0_001_10011100;
	12'b0_000_10100000 : r_w_inv <= 12'b0_001_10011010;
	12'b0_000_10100001 : r_w_inv <= 12'b0_001_10011000;
	12'b0_000_10100010 : r_w_inv <= 12'b0_001_10010101;
	12'b0_000_10100011 : r_w_inv <= 12'b0_001_10010011;
	12'b0_000_10100100 : r_w_inv <= 12'b0_001_10010000;
	12'b0_000_10100101 : r_w_inv <= 12'b0_001_10001110;
	12'b0_000_10100110 : r_w_inv <= 12'b0_001_10001011;
	12'b0_000_10100111 : r_w_inv <= 12'b0_001_10001001;
	12'b0_000_10101000 : r_w_inv <= 12'b0_001_10000110;
	12'b0_000_10101001 : r_w_inv <= 12'b0_001_10000100;
	12'b0_000_10101010 : r_w_inv <= 12'b0_001_10000010;
	12'b0_000_10101011 : r_w_inv <= 12'b0_001_01111111;
	12'b0_000_10101100 : r_w_inv <= 12'b0_001_01111110;
	12'b0_000_10101101 : r_w_inv <= 12'b0_001_01111011;
	12'b0_000_10101110 : r_w_inv <= 12'b0_001_01111001;
	12'b0_000_10101111 : r_w_inv <= 12'b0_001_01110111;
	12'b0_000_10110000 : r_w_inv <= 12'b0_001_01110101;
	12'b0_000_10110001 : r_w_inv <= 12'b0_001_01110010;
	12'b0_000_10110010 : r_w_inv <= 12'b0_001_01110000;
	12'b0_000_10110011 : r_w_inv <= 12'b0_001_01101110;
	12'b0_000_10110100 : r_w_inv <= 12'b0_001_01101100;
	12'b0_000_10110101 : r_w_inv <= 12'b0_001_01101010;
	12'b0_000_10110110 : r_w_inv <= 12'b0_001_01101001;
	12'b0_000_10110111 : r_w_inv <= 12'b0_001_01100111;
	12'b0_000_10111000 : r_w_inv <= 12'b0_001_01100101;
	12'b0_000_10111001 : r_w_inv <= 12'b0_001_01100011;
	12'b0_000_10111010 : r_w_inv <= 12'b0_001_01100001;
	12'b0_000_10111011 : r_w_inv <= 12'b0_001_01011111;
	12'b0_000_10111100 : r_w_inv <= 12'b0_001_01011101;
	12'b0_000_10111101 : r_w_inv <= 12'b0_001_01011011;
	12'b0_000_10111110 : r_w_inv <= 12'b0_001_01011001;
	12'b0_000_10111111 : r_w_inv <= 12'b0_001_01010111;
	12'b0_000_11000000 : r_w_inv <= 12'b0_001_01010101;
	12'b0_000_11000001 : r_w_inv <= 12'b0_001_01010100;
	12'b0_000_11000010 : r_w_inv <= 12'b0_001_01010010;
	12'b0_000_11000011 : r_w_inv <= 12'b0_001_01010000;
	12'b0_000_11000100 : r_w_inv <= 12'b0_001_01001111;
	12'b0_000_11000101 : r_w_inv <= 12'b0_001_01001101;
	12'b0_000_11000110 : r_w_inv <= 12'b0_001_01001011;
	12'b0_000_11000111 : r_w_inv <= 12'b0_001_01001001;
	12'b0_000_11001000 : r_w_inv <= 12'b0_001_01001000;
	12'b0_000_11001001 : r_w_inv <= 12'b0_001_01000110;
	12'b0_000_11001010 : r_w_inv <= 12'b0_001_01000100;
	12'b0_000_11001011 : r_w_inv <= 12'b0_001_01000011;
	12'b0_000_11001100 : r_w_inv <= 12'b0_001_01000010;
	12'b0_000_11001101 : r_w_inv <= 12'b0_001_01000000;
	12'b0_000_11001110 : r_w_inv <= 12'b0_001_00111110;
	12'b0_000_11001111 : r_w_inv <= 12'b0_001_00111101;
	12'b0_000_11010000 : r_w_inv <= 12'b0_001_00111011;
	12'b0_000_11010001 : r_w_inv <= 12'b0_001_00111010;
	12'b0_000_11010010 : r_w_inv <= 12'b0_001_00111000;
	12'b0_000_11010011 : r_w_inv <= 12'b0_001_00110111;
	12'b0_000_11010100 : r_w_inv <= 12'b0_001_00110101;
	12'b0_000_11010101 : r_w_inv <= 12'b0_001_00110100;
	12'b0_000_11010110 : r_w_inv <= 12'b0_001_00110011;
	12'b0_000_11010111 : r_w_inv <= 12'b0_001_00110001;
	12'b0_000_11011000 : r_w_inv <= 12'b0_001_00110000;
	12'b0_000_11011001 : r_w_inv <= 12'b0_001_00101110;
	12'b0_000_11011010 : r_w_inv <= 12'b0_001_00101101;
	12'b0_000_11011011 : r_w_inv <= 12'b0_001_00101011;
	12'b0_000_11011100 : r_w_inv <= 12'b0_001_00101010;
	12'b0_000_11011101 : r_w_inv <= 12'b0_001_00101001;
	12'b0_000_11011110 : r_w_inv <= 12'b0_001_00100111;
	12'b0_000_11011111 : r_w_inv <= 12'b0_001_00100110;
	12'b0_000_11100000 : r_w_inv <= 12'b0_001_00100101;
	12'b0_000_11100001 : r_w_inv <= 12'b0_001_00100100;
	12'b0_000_11100010 : r_w_inv <= 12'b0_001_00100010;
	12'b0_000_11100011 : r_w_inv <= 12'b0_001_00100001;
	12'b0_000_11100100 : r_w_inv <= 12'b0_001_00100000;
	12'b0_000_11100101 : r_w_inv <= 12'b0_001_00011110;
	12'b0_000_11100110 : r_w_inv <= 12'b0_001_00011101;
	12'b0_000_11100111 : r_w_inv <= 12'b0_001_00011100;
	12'b0_000_11101000 : r_w_inv <= 12'b0_001_00011011;
	12'b0_000_11101001 : r_w_inv <= 12'b0_001_00011001;
	12'b0_000_11101010 : r_w_inv <= 12'b0_001_00011000;
	12'b0_000_11101011 : r_w_inv <= 12'b0_001_00010111;
	12'b0_000_11101100 : r_w_inv <= 12'b0_001_00010110;
	12'b0_000_11101101 : r_w_inv <= 12'b0_001_00010101;
	12'b0_000_11101110 : r_w_inv <= 12'b0_001_00010100;
	12'b0_000_11101111 : r_w_inv <= 12'b0_001_00010010;
	12'b0_000_11110000 : r_w_inv <= 12'b0_001_00010001;
	12'b0_000_11110001 : r_w_inv <= 12'b0_001_00010000;
	12'b0_000_11110010 : r_w_inv <= 12'b0_001_00001111;
	12'b0_000_11110011 : r_w_inv <= 12'b0_001_00001110;
	12'b0_000_11110100 : r_w_inv <= 12'b0_001_00001101;
	12'b0_000_11110101 : r_w_inv <= 12'b0_001_00001100;
	12'b0_000_11110110 : r_w_inv <= 12'b0_001_00001011;
	12'b0_000_11110111 : r_w_inv <= 12'b0_001_00001010;
	12'b0_000_11111000 : r_w_inv <= 12'b0_001_00001000;
	12'b0_000_11111001 : r_w_inv <= 12'b0_001_00000111;
	12'b0_000_11111010 : r_w_inv <= 12'b0_001_00000110;
	12'b0_000_11111011 : r_w_inv <= 12'b0_001_00000101;
	12'b0_000_11111100 : r_w_inv <= 12'b0_001_00000100;
	12'b0_000_11111101 : r_w_inv <= 12'b0_001_00000011;
	12'b0_000_11111110 : r_w_inv <= 12'b0_001_00000010;
	12'b0_000_11111111 : r_w_inv <= 12'b0_001_00000001;
	12'b0_001_00000000 : r_w_inv <= 12'b0_001_00000000;
	12'b0_001_00000001 : r_w_inv <= 12'b0_000_11111111;
	12'b0_001_00000010 : r_w_inv <= 12'b0_000_11111110;
	12'b0_001_00000011 : r_w_inv <= 12'b0_000_11111101;
	12'b0_001_00000100 : r_w_inv <= 12'b0_000_11111100;
	12'b0_001_00000101 : r_w_inv <= 12'b0_000_11111011;
	12'b0_001_00000110 : r_w_inv <= 12'b0_000_11111010;
	12'b0_001_00000111 : r_w_inv <= 12'b0_000_11111001;
	12'b0_001_00001000 : r_w_inv <= 12'b0_000_11111000;
	12'b0_001_00001001 : r_w_inv <= 12'b0_000_11110111;
	12'b0_001_00001010 : r_w_inv <= 12'b0_000_11110110;
	12'b0_001_00001011 : r_w_inv <= 12'b0_000_11110101;
	12'b0_001_00001100 : r_w_inv <= 12'b0_000_11110101;
	12'b0_001_00001101 : r_w_inv <= 12'b0_000_11110100;
	12'b0_001_00001110 : r_w_inv <= 12'b0_000_11110011;
	12'b0_001_00001111 : r_w_inv <= 12'b0_000_11110010;
	12'b0_001_00010000 : r_w_inv <= 12'b0_000_11110001;
	12'b0_001_00010001 : r_w_inv <= 12'b0_000_11110000;
	12'b0_001_00010010 : r_w_inv <= 12'b0_000_11101111;
	12'b0_001_00010011 : r_w_inv <= 12'b0_000_11101110;
	12'b0_001_00010100 : r_w_inv <= 12'b0_000_11101101;
	12'b0_001_00010101 : r_w_inv <= 12'b0_000_11101101;
	12'b0_001_00010110 : r_w_inv <= 12'b0_000_11101100;
	12'b0_001_00010111 : r_w_inv <= 12'b0_000_11101011;
	12'b0_001_00011000 : r_w_inv <= 12'b0_000_11101010;
	12'b0_001_00011001 : r_w_inv <= 12'b0_000_11101001;
	12'b0_001_00011010 : r_w_inv <= 12'b0_000_11101001;
	12'b0_001_00011011 : r_w_inv <= 12'b0_000_11101000;
	12'b0_001_00011100 : r_w_inv <= 12'b0_000_11100111;
	12'b0_001_00011101 : r_w_inv <= 12'b0_000_11100110;
	12'b0_001_00011110 : r_w_inv <= 12'b0_000_11100101;
	12'b0_001_00011111 : r_w_inv <= 12'b0_000_11100100;
	12'b0_001_00100000 : r_w_inv <= 12'b0_000_11100100;
	12'b0_001_00100001 : r_w_inv <= 12'b0_000_11100011;
	12'b0_001_00100010 : r_w_inv <= 12'b0_000_11100010;
	12'b0_001_00100011 : r_w_inv <= 12'b0_000_11100001;
	12'b0_001_00100100 : r_w_inv <= 12'b0_000_11100001;
	12'b0_001_00100101 : r_w_inv <= 12'b0_000_11100000;
	12'b0_001_00100110 : r_w_inv <= 12'b0_000_11011111;
	12'b0_001_00100111 : r_w_inv <= 12'b0_000_11011110;
	12'b0_001_00101000 : r_w_inv <= 12'b0_000_11011101;
	12'b0_001_00101001 : r_w_inv <= 12'b0_000_11011101;
	12'b0_001_00101010 : r_w_inv <= 12'b0_000_11011100;
	12'b0_001_00101011 : r_w_inv <= 12'b0_000_11011011;
	12'b0_001_00101100 : r_w_inv <= 12'b0_000_11011011;
	12'b0_001_00101101 : r_w_inv <= 12'b0_000_11011010;
	12'b0_001_00101110 : r_w_inv <= 12'b0_000_11011001;
	12'b0_001_00101111 : r_w_inv <= 12'b0_000_11011000;
	12'b0_001_00110000 : r_w_inv <= 12'b0_000_11011000;
	12'b0_001_00110001 : r_w_inv <= 12'b0_000_11010111;
	12'b0_001_00110010 : r_w_inv <= 12'b0_000_11010110;
	12'b0_001_00110011 : r_w_inv <= 12'b0_000_11010110;
	12'b0_001_00110100 : r_w_inv <= 12'b0_000_11010101;
	12'b0_001_00110101 : r_w_inv <= 12'b0_000_11010100;
	12'b0_001_00110110 : r_w_inv <= 12'b0_000_11010100;
	12'b0_001_00110111 : r_w_inv <= 12'b0_000_11010011;
	12'b0_001_00111000 : r_w_inv <= 12'b0_000_11010010;
	12'b0_001_00111001 : r_w_inv <= 12'b0_000_11010001;
	12'b0_001_00111010 : r_w_inv <= 12'b0_000_11010001;
	12'b0_001_00111011 : r_w_inv <= 12'b0_000_11010000;
	12'b0_001_00111100 : r_w_inv <= 12'b0_000_11001111;
	12'b0_001_00111101 : r_w_inv <= 12'b0_000_11001111;
	12'b0_001_00111110 : r_w_inv <= 12'b0_000_11001110;
	12'b0_001_00111111 : r_w_inv <= 12'b0_000_11001101;
	12'b0_001_01000000 : r_w_inv <= 12'b0_000_11001101;
	12'b0_001_01000001 : r_w_inv <= 12'b0_000_11001100;
	12'b0_001_01000010 : r_w_inv <= 12'b0_000_11001100;
	12'b0_001_01000011 : r_w_inv <= 12'b0_000_11001011;
	12'b0_001_01000100 : r_w_inv <= 12'b0_000_11001010;
	12'b0_001_01000101 : r_w_inv <= 12'b0_000_11001010;
	12'b0_001_01000110 : r_w_inv <= 12'b0_000_11001001;
	12'b0_001_01000111 : r_w_inv <= 12'b0_000_11001000;
	12'b0_001_01001000 : r_w_inv <= 12'b0_000_11001000;
	12'b0_001_01001001 : r_w_inv <= 12'b0_000_11000111;
	12'b0_001_01001010 : r_w_inv <= 12'b0_000_11000111;
	12'b0_001_01001011 : r_w_inv <= 12'b0_000_11000110;
	12'b0_001_01001100 : r_w_inv <= 12'b0_000_11000110;
	12'b0_001_01001101 : r_w_inv <= 12'b0_000_11000101;
	12'b0_001_01001110 : r_w_inv <= 12'b0_000_11000100;
	12'b0_001_01001111 : r_w_inv <= 12'b0_000_11000100;
	12'b0_001_01010000 : r_w_inv <= 12'b0_000_11000011;
	12'b0_001_01010001 : r_w_inv <= 12'b0_000_11000011;
	12'b0_001_01010010 : r_w_inv <= 12'b0_000_11000010;
	12'b0_001_01010011 : r_w_inv <= 12'b0_000_11000001;
	12'b0_001_01010100 : r_w_inv <= 12'b0_000_11000001;
	12'b0_001_01010101 : r_w_inv <= 12'b0_000_11000000;
	12'b0_001_01010110 : r_w_inv <= 12'b0_000_11000000;
	12'b0_001_01010111 : r_w_inv <= 12'b0_000_10111111;
	12'b0_001_01011000 : r_w_inv <= 12'b0_000_10111111;
	12'b0_001_01011001 : r_w_inv <= 12'b0_000_10111110;
	12'b0_001_01011010 : r_w_inv <= 12'b0_000_10111101;
	12'b0_001_01011011 : r_w_inv <= 12'b0_000_10111101;
	12'b0_001_01011100 : r_w_inv <= 12'b0_000_10111100;
	12'b0_001_01011101 : r_w_inv <= 12'b0_000_10111100;
	12'b0_001_01011110 : r_w_inv <= 12'b0_000_10111011;
	12'b0_001_01011111 : r_w_inv <= 12'b0_000_10111011;
	12'b0_001_01100000 : r_w_inv <= 12'b0_000_10111010;
	12'b0_001_01100001 : r_w_inv <= 12'b0_000_10111010;
	12'b0_001_01100010 : r_w_inv <= 12'b0_000_10111001;
	12'b0_001_01100011 : r_w_inv <= 12'b0_000_10111001;
	12'b0_001_01100100 : r_w_inv <= 12'b0_000_10111000;
	12'b0_001_01100101 : r_w_inv <= 12'b0_000_10111000;
	12'b0_001_01100110 : r_w_inv <= 12'b0_000_10110111;
	12'b0_001_01100111 : r_w_inv <= 12'b0_000_10110111;
	12'b0_001_01101000 : r_w_inv <= 12'b0_000_10110110;
	12'b0_001_01101001 : r_w_inv <= 12'b0_000_10110110;
	12'b0_001_01101010 : r_w_inv <= 12'b0_000_10110101;
	12'b0_001_01101011 : r_w_inv <= 12'b0_000_10110101;
	12'b0_001_01101100 : r_w_inv <= 12'b0_000_10110100;
	12'b0_001_01101101 : r_w_inv <= 12'b0_000_10110100;
	12'b0_001_01101110 : r_w_inv <= 12'b0_000_10110011;
	12'b0_001_01101111 : r_w_inv <= 12'b0_000_10110011;
	12'b0_001_01110000 : r_w_inv <= 12'b0_000_10110010;
	12'b0_001_01110001 : r_w_inv <= 12'b0_000_10110010;
	12'b0_001_01110010 : r_w_inv <= 12'b0_000_10110001;
	12'b0_001_01110011 : r_w_inv <= 12'b0_000_10110001;
	12'b0_001_01110100 : r_w_inv <= 12'b0_000_10110000;
	12'b0_001_01110101 : r_w_inv <= 12'b0_000_10110000;
	12'b0_001_01110110 : r_w_inv <= 12'b0_000_10101111;
	12'b0_001_01110111 : r_w_inv <= 12'b0_000_10101111;
	12'b0_001_01111000 : r_w_inv <= 12'b0_000_10101110;
	12'b0_001_01111001 : r_w_inv <= 12'b0_000_10101110;
	12'b0_001_01111010 : r_w_inv <= 12'b0_000_10101101;
	12'b0_001_01111011 : r_w_inv <= 12'b0_000_10101101;
	12'b0_001_01111100 : r_w_inv <= 12'b0_000_10101101;
	12'b0_001_01111101 : r_w_inv <= 12'b0_000_10101100;
	12'b0_001_01111110 : r_w_inv <= 12'b0_000_10101100;
	12'b0_001_01111111 : r_w_inv <= 12'b0_000_10101011;
	12'b0_001_10000000 : r_w_inv <= 12'b0_000_10101011;
	12'b0_001_10000001 : r_w_inv <= 12'b0_000_10101010;
	12'b0_001_10000010 : r_w_inv <= 12'b0_000_10101010;
	12'b0_001_10000011 : r_w_inv <= 12'b0_000_10101001;
	12'b0_001_10000100 : r_w_inv <= 12'b0_000_10101001;
	12'b0_001_10000101 : r_w_inv <= 12'b0_000_10101001;
	12'b0_001_10000110 : r_w_inv <= 12'b0_000_10101000;
	12'b0_001_10000111 : r_w_inv <= 12'b0_000_10101000;
	12'b0_001_10001000 : r_w_inv <= 12'b0_000_10100111;
	12'b0_001_10001001 : r_w_inv <= 12'b0_000_10100111;
	12'b0_001_10001010 : r_w_inv <= 12'b0_000_10100110;
	12'b0_001_10001011 : r_w_inv <= 12'b0_000_10100110;
	12'b0_001_10001100 : r_w_inv <= 12'b0_000_10100110;
	12'b0_001_10001101 : r_w_inv <= 12'b0_000_10100101;
	12'b0_001_10001110 : r_w_inv <= 12'b0_000_10100101;
	12'b0_001_10001111 : r_w_inv <= 12'b0_000_10100100;
	12'b0_001_10010000 : r_w_inv <= 12'b0_000_10100100;
	12'b0_001_10010001 : r_w_inv <= 12'b0_000_10100011;
	12'b0_001_10010010 : r_w_inv <= 12'b0_000_10100011;
	12'b0_001_10010011 : r_w_inv <= 12'b0_000_10100011;
	12'b0_001_10010100 : r_w_inv <= 12'b0_000_10100010;
	12'b0_001_10010101 : r_w_inv <= 12'b0_000_10100010;
	12'b0_001_10010110 : r_w_inv <= 12'b0_000_10100010;
	12'b0_001_10010111 : r_w_inv <= 12'b0_000_10100001;
	12'b0_001_10011000 : r_w_inv <= 12'b0_000_10100001;
	12'b0_001_10011001 : r_w_inv <= 12'b0_000_10100000;
	12'b0_001_10011010 : r_w_inv <= 12'b0_000_10100000;
	12'b0_001_10011011 : r_w_inv <= 12'b0_000_10100000;
	12'b0_001_10011100 : r_w_inv <= 12'b0_000_10011111;
	12'b0_001_10011101 : r_w_inv <= 12'b0_000_10011111;
	12'b0_001_10011110 : r_w_inv <= 12'b0_000_10011110;
	12'b0_001_10011111 : r_w_inv <= 12'b0_000_10011110;
	12'b0_001_10100000 : r_w_inv <= 12'b0_000_10011110;
	12'b0_001_10100001 : r_w_inv <= 12'b0_000_10011101;
	12'b0_001_10100010 : r_w_inv <= 12'b0_000_10011101;
	12'b0_001_10100011 : r_w_inv <= 12'b0_000_10011100;
	12'b0_001_10100100 : r_w_inv <= 12'b0_000_10011100;
	12'b0_001_10100101 : r_w_inv <= 12'b0_000_10011100;
	12'b0_001_10100110 : r_w_inv <= 12'b0_000_10011011;
	12'b0_001_10100111 : r_w_inv <= 12'b0_000_10011011;
	12'b0_001_10101000 : r_w_inv <= 12'b0_000_10011011;
	12'b0_001_10101001 : r_w_inv <= 12'b0_000_10011010;
	12'b0_001_10101010 : r_w_inv <= 12'b0_000_10011010;
	12'b0_001_10101011 : r_w_inv <= 12'b0_000_10011001;
	12'b0_001_10101100 : r_w_inv <= 12'b0_000_10011001;
	12'b0_001_10101101 : r_w_inv <= 12'b0_000_10011001;
	12'b0_001_10101110 : r_w_inv <= 12'b0_000_10011000;
	12'b0_001_10101111 : r_w_inv <= 12'b0_000_10011000;
	12'b0_001_10110000 : r_w_inv <= 12'b0_000_10011000;
	12'b0_001_10110001 : r_w_inv <= 12'b0_000_10010111;
	12'b0_001_10110010 : r_w_inv <= 12'b0_000_10010111;
	12'b0_001_10110011 : r_w_inv <= 12'b0_000_10010111;
	12'b0_001_10110100 : r_w_inv <= 12'b0_000_10010110;
	12'b0_001_10110101 : r_w_inv <= 12'b0_000_10010110;
	12'b0_001_10110110 : r_w_inv <= 12'b0_000_10010110;
	12'b0_001_10110111 : r_w_inv <= 12'b0_000_10010101;
	12'b0_001_10111000 : r_w_inv <= 12'b0_000_10010101;
	12'b0_001_10111001 : r_w_inv <= 12'b0_000_10010101;
	12'b0_001_10111010 : r_w_inv <= 12'b0_000_10010100;
	12'b0_001_10111011 : r_w_inv <= 12'b0_000_10010100;
	12'b0_001_10111100 : r_w_inv <= 12'b0_000_10010100;
	12'b0_001_10111101 : r_w_inv <= 12'b0_000_10010011;
	12'b0_001_10111110 : r_w_inv <= 12'b0_000_10010011;
	12'b0_001_10111111 : r_w_inv <= 12'b0_000_10010011;
	12'b0_001_11000000 : r_w_inv <= 12'b0_000_10010010;
	12'b0_001_11000001 : r_w_inv <= 12'b0_000_10010010;
	12'b0_001_11000010 : r_w_inv <= 12'b0_000_10010010;
	12'b0_001_11000011 : r_w_inv <= 12'b0_000_10010001;
	12'b0_001_11000100 : r_w_inv <= 12'b0_000_10010001;
	12'b0_001_11000101 : r_w_inv <= 12'b0_000_10010001;
	12'b0_001_11000110 : r_w_inv <= 12'b0_000_10010000;
	12'b0_001_11000111 : r_w_inv <= 12'b0_000_10010000;
	12'b0_001_11001000 : r_w_inv <= 12'b0_000_10010000;
	12'b0_001_11001001 : r_w_inv <= 12'b0_000_10001111;
	12'b0_001_11001010 : r_w_inv <= 12'b0_000_10001111;
	12'b0_001_11001011 : r_w_inv <= 12'b0_000_10001111;
	12'b0_001_11001100 : r_w_inv <= 12'b0_000_10001111;
	12'b0_001_11001101 : r_w_inv <= 12'b0_000_10001110;
	12'b0_001_11001110 : r_w_inv <= 12'b0_000_10001110;
	12'b0_001_11001111 : r_w_inv <= 12'b0_000_10001110;
	12'b0_001_11010000 : r_w_inv <= 12'b0_000_10001101;
	12'b0_001_11010001 : r_w_inv <= 12'b0_000_10001101;
	12'b0_001_11010010 : r_w_inv <= 12'b0_000_10001101;
	12'b0_001_11010011 : r_w_inv <= 12'b0_000_10001100;
	12'b0_001_11010100 : r_w_inv <= 12'b0_000_10001100;
	12'b0_001_11010101 : r_w_inv <= 12'b0_000_10001100;
	12'b0_001_11010110 : r_w_inv <= 12'b0_000_10001100;
	12'b0_001_11010111 : r_w_inv <= 12'b0_000_10001011;
	12'b0_001_11011000 : r_w_inv <= 12'b0_000_10001011;
	12'b0_001_11011001 : r_w_inv <= 12'b0_000_10001011;
	12'b0_001_11011010 : r_w_inv <= 12'b0_000_10001010;
	12'b0_001_11011011 : r_w_inv <= 12'b0_000_10001010;
	12'b0_001_11011100 : r_w_inv <= 12'b0_000_10001010;
	12'b0_001_11011101 : r_w_inv <= 12'b0_000_10001001;
	12'b0_001_11011110 : r_w_inv <= 12'b0_000_10001001;
	12'b0_001_11011111 : r_w_inv <= 12'b0_000_10001001;
	12'b0_001_11100000 : r_w_inv <= 12'b0_000_10001001;
	12'b0_001_11100001 : r_w_inv <= 12'b0_000_10001000;
	12'b0_001_11100010 : r_w_inv <= 12'b0_000_10001000;
	12'b0_001_11100011 : r_w_inv <= 12'b0_000_10001000;
	12'b0_001_11100100 : r_w_inv <= 12'b0_000_10000111;
	12'b0_001_11100101 : r_w_inv <= 12'b0_000_10000111;
	12'b0_001_11100110 : r_w_inv <= 12'b0_000_10000111;
	12'b0_001_11100111 : r_w_inv <= 12'b0_000_10000111;
	12'b0_001_11101000 : r_w_inv <= 12'b0_000_10000110;
	12'b0_001_11101001 : r_w_inv <= 12'b0_000_10000110;
	12'b0_001_11101010 : r_w_inv <= 12'b0_000_10000110;
	12'b0_001_11101011 : r_w_inv <= 12'b0_000_10000101;
	12'b0_001_11101100 : r_w_inv <= 12'b0_000_10000101;
	12'b0_001_11101101 : r_w_inv <= 12'b0_000_10000101;
	12'b0_001_11101110 : r_w_inv <= 12'b0_000_10000101;
	12'b0_001_11101111 : r_w_inv <= 12'b0_000_10000100;
	12'b0_001_11110000 : r_w_inv <= 12'b0_000_10000100;
	12'b0_001_11110001 : r_w_inv <= 12'b0_000_10000100;
	12'b0_001_11110010 : r_w_inv <= 12'b0_000_10000100;
	12'b0_001_11110011 : r_w_inv <= 12'b0_000_10000011;
	12'b0_001_11110100 : r_w_inv <= 12'b0_000_10000011;
	12'b0_001_11110101 : r_w_inv <= 12'b0_000_10000011;
	12'b0_001_11110110 : r_w_inv <= 12'b0_000_10000011;
	12'b0_001_11110111 : r_w_inv <= 12'b0_000_10000010;
	12'b0_001_11111000 : r_w_inv <= 12'b0_000_10000010;
	12'b0_001_11111001 : r_w_inv <= 12'b0_000_10000010;
	12'b0_001_11111010 : r_w_inv <= 12'b0_000_10000010;
	12'b0_001_11111011 : r_w_inv <= 12'b0_000_10000001;
	12'b0_001_11111100 : r_w_inv <= 12'b0_000_10000001;
	12'b0_001_11111101 : r_w_inv <= 12'b0_000_10000001;
	12'b0_001_11111110 : r_w_inv <= 12'b0_000_10000001;
	12'b0_001_11111111 : r_w_inv <= 12'b0_000_10000000;
	12'b0_010_00000000 : r_w_inv <= 12'b0_000_10000000;
	12'b0_010_00000001 : r_w_inv <= 12'b0_000_10000000;
	12'b0_010_00000010 : r_w_inv <= 12'b0_000_10000000;
	12'b0_010_00000011 : r_w_inv <= 12'b0_000_01111111;
	12'b0_010_00000100 : r_w_inv <= 12'b0_000_01111111;
	12'b0_010_00000101 : r_w_inv <= 12'b0_000_01111111;
	12'b0_010_00000110 : r_w_inv <= 12'b0_000_01111111;
	12'b0_010_00000111 : r_w_inv <= 12'b0_000_01111110;
	12'b0_010_00001000 : r_w_inv <= 12'b0_000_01111110;
	12'b0_010_00001001 : r_w_inv <= 12'b0_000_01111110;
	12'b0_010_00001010 : r_w_inv <= 12'b0_000_01111110;
	12'b0_010_00001011 : r_w_inv <= 12'b0_000_01111101;
	12'b0_010_00001100 : r_w_inv <= 12'b0_000_01111101;
	12'b0_010_00001101 : r_w_inv <= 12'b0_000_01111101;
	12'b0_010_00001110 : r_w_inv <= 12'b0_000_01111101;
	12'b0_010_00001111 : r_w_inv <= 12'b0_000_01111100;
	12'b0_010_00010000 : r_w_inv <= 12'b0_000_01111100;
	12'b0_010_00010001 : r_w_inv <= 12'b0_000_01111100;
	12'b0_010_00010010 : r_w_inv <= 12'b0_000_01111100;
	12'b0_010_00010011 : r_w_inv <= 12'b0_000_01111011;
	12'b0_010_00010100 : r_w_inv <= 12'b0_000_01111011;
	12'b0_010_00010101 : r_w_inv <= 12'b0_000_01111011;
	12'b0_010_00010110 : r_w_inv <= 12'b0_000_01111011;
	12'b0_010_00010111 : r_w_inv <= 12'b0_000_01111011;
	12'b0_010_00011000 : r_w_inv <= 12'b0_000_01111010;
	12'b0_010_00011001 : r_w_inv <= 12'b0_000_01111010;
	12'b0_010_00011010 : r_w_inv <= 12'b0_000_01111010;
	12'b0_010_00011011 : r_w_inv <= 12'b0_000_01111010;
	12'b0_010_00011100 : r_w_inv <= 12'b0_000_01111001;
	12'b0_010_00011101 : r_w_inv <= 12'b0_000_01111001;
	12'b0_010_00011110 : r_w_inv <= 12'b0_000_01111001;
	12'b0_010_00011111 : r_w_inv <= 12'b0_000_01111001;
	12'b0_010_00100000 : r_w_inv <= 12'b0_000_01111000;
	12'b0_010_00100001 : r_w_inv <= 12'b0_000_01111000;
	12'b0_010_00100010 : r_w_inv <= 12'b0_000_01111000;
	12'b0_010_00100011 : r_w_inv <= 12'b0_000_01111000;
	12'b0_010_00100100 : r_w_inv <= 12'b0_000_01111000;
	12'b0_010_00100101 : r_w_inv <= 12'b0_000_01110111;
	12'b0_010_00100110 : r_w_inv <= 12'b0_000_01110111;
	12'b0_010_00100111 : r_w_inv <= 12'b0_000_01110111;
	12'b0_010_00101000 : r_w_inv <= 12'b0_000_01110111;
	12'b0_010_00101001 : r_w_inv <= 12'b0_000_01110111;
	12'b0_010_00101010 : r_w_inv <= 12'b0_000_01110110;
	12'b0_010_00101011 : r_w_inv <= 12'b0_000_01110110;
	12'b0_010_00101100 : r_w_inv <= 12'b0_000_01110110;
	12'b0_010_00101101 : r_w_inv <= 12'b0_000_01110110;
	12'b0_010_00101110 : r_w_inv <= 12'b0_000_01110101;
	12'b0_010_00101111 : r_w_inv <= 12'b0_000_01110101;
	12'b0_010_00110000 : r_w_inv <= 12'b0_000_01110101;
	12'b0_010_00110001 : r_w_inv <= 12'b0_000_01110101;
	12'b0_010_00110010 : r_w_inv <= 12'b0_000_01110101;
	12'b0_010_00110011 : r_w_inv <= 12'b0_000_01110100;
	12'b0_010_00110100 : r_w_inv <= 12'b0_000_01110100;
	12'b0_010_00110101 : r_w_inv <= 12'b0_000_01110100;
	12'b0_010_00110110 : r_w_inv <= 12'b0_000_01110100;
	12'b0_010_00110111 : r_w_inv <= 12'b0_000_01110100;
	12'b0_010_00111000 : r_w_inv <= 12'b0_000_01110011;
	12'b0_010_00111001 : r_w_inv <= 12'b0_000_01110011;
	12'b0_010_00111010 : r_w_inv <= 12'b0_000_01110011;
	12'b0_010_00111011 : r_w_inv <= 12'b0_000_01110011;
	12'b0_010_00111100 : r_w_inv <= 12'b0_000_01110011;
	12'b0_010_00111101 : r_w_inv <= 12'b0_000_01110010;
	12'b0_010_00111110 : r_w_inv <= 12'b0_000_01110010;
	12'b0_010_00111111 : r_w_inv <= 12'b0_000_01110010;
	12'b0_010_01000000 : r_w_inv <= 12'b0_000_01110010;
	12'b0_010_01000001 : r_w_inv <= 12'b0_000_01110010;
	12'b0_010_01000010 : r_w_inv <= 12'b0_000_01110001;
	12'b0_010_01000011 : r_w_inv <= 12'b0_000_01110001;
	12'b0_010_01000100 : r_w_inv <= 12'b0_000_01110001;
	12'b0_010_01000101 : r_w_inv <= 12'b0_000_01110001;
	12'b0_010_01000110 : r_w_inv <= 12'b0_000_01110001;
	12'b0_010_01000111 : r_w_inv <= 12'b0_000_01110000;
	12'b0_010_01001000 : r_w_inv <= 12'b0_000_01110000;
	12'b0_010_01001001 : r_w_inv <= 12'b0_000_01110000;
	12'b0_010_01001010 : r_w_inv <= 12'b0_000_01110000;
	12'b0_010_01001011 : r_w_inv <= 12'b0_000_01110000;
	12'b0_010_01001100 : r_w_inv <= 12'b0_000_01101111;
	12'b0_010_01001101 : r_w_inv <= 12'b0_000_01101111;
	12'b0_010_01001110 : r_w_inv <= 12'b0_000_01101111;
	12'b0_010_01001111 : r_w_inv <= 12'b0_000_01101111;
	12'b0_010_01010000 : r_w_inv <= 12'b0_000_01101111;
	12'b0_010_01010001 : r_w_inv <= 12'b0_000_01101111;
	12'b0_010_01010010 : r_w_inv <= 12'b0_000_01101110;
	12'b0_010_01010011 : r_w_inv <= 12'b0_000_01101110;
	12'b0_010_01010100 : r_w_inv <= 12'b0_000_01101110;
	12'b0_010_01010101 : r_w_inv <= 12'b0_000_01101110;
	12'b0_010_01010110 : r_w_inv <= 12'b0_000_01101110;
	12'b0_010_01010111 : r_w_inv <= 12'b0_000_01101101;
	12'b0_010_01011000 : r_w_inv <= 12'b0_000_01101101;
	12'b0_010_01011001 : r_w_inv <= 12'b0_000_01101101;
	12'b0_010_01011010 : r_w_inv <= 12'b0_000_01101101;
	12'b0_010_01011011 : r_w_inv <= 12'b0_000_01101101;
	12'b0_010_01011100 : r_w_inv <= 12'b0_000_01101101;
	12'b0_010_01011101 : r_w_inv <= 12'b0_000_01101100;
	12'b0_010_01011110 : r_w_inv <= 12'b0_000_01101100;
	12'b0_010_01011111 : r_w_inv <= 12'b0_000_01101100;
	12'b0_010_01100000 : r_w_inv <= 12'b0_000_01101100;
	12'b0_010_01100001 : r_w_inv <= 12'b0_000_01101100;
	12'b0_010_01100010 : r_w_inv <= 12'b0_000_01101011;
	12'b0_010_01100011 : r_w_inv <= 12'b0_000_01101011;
	12'b0_010_01100100 : r_w_inv <= 12'b0_000_01101011;
	12'b0_010_01100101 : r_w_inv <= 12'b0_000_01101011;
	12'b0_010_01100110 : r_w_inv <= 12'b0_000_01101011;
	12'b0_010_01100111 : r_w_inv <= 12'b0_000_01101011;
	12'b0_010_01101000 : r_w_inv <= 12'b0_000_01101010;
	12'b0_010_01101001 : r_w_inv <= 12'b0_000_01101010;
	12'b0_010_01101010 : r_w_inv <= 12'b0_000_01101010;
	12'b0_010_01101011 : r_w_inv <= 12'b0_000_01101010;
	12'b0_010_01101100 : r_w_inv <= 12'b0_000_01101010;
	12'b0_010_01101101 : r_w_inv <= 12'b0_000_01101010;
	12'b0_010_01101110 : r_w_inv <= 12'b0_000_01101001;
	12'b0_010_01101111 : r_w_inv <= 12'b0_000_01101001;
	12'b0_010_01110000 : r_w_inv <= 12'b0_000_01101001;
	12'b0_010_01110001 : r_w_inv <= 12'b0_000_01101001;
	12'b0_010_01110010 : r_w_inv <= 12'b0_000_01101001;
	12'b0_010_01110011 : r_w_inv <= 12'b0_000_01101001;
	12'b0_010_01110100 : r_w_inv <= 12'b0_000_01101000;
	12'b0_010_01110101 : r_w_inv <= 12'b0_000_01101000;
	12'b0_010_01110110 : r_w_inv <= 12'b0_000_01101000;
	12'b0_010_01110111 : r_w_inv <= 12'b0_000_01101000;
	12'b0_010_01111000 : r_w_inv <= 12'b0_000_01101000;
	12'b0_010_01111001 : r_w_inv <= 12'b0_000_01101000;
	12'b0_010_01111010 : r_w_inv <= 12'b0_000_01100111;
	12'b0_010_01111011 : r_w_inv <= 12'b0_000_01100111;
	12'b0_010_01111100 : r_w_inv <= 12'b0_000_01100111;
	12'b0_010_01111101 : r_w_inv <= 12'b0_000_01100111;
	12'b0_010_01111110 : r_w_inv <= 12'b0_000_01100111;
	12'b0_010_01111111 : r_w_inv <= 12'b0_000_01100111;
	12'b0_010_10000000 : r_w_inv <= 12'b0_000_01100110;
	12'b0_010_10000001 : r_w_inv <= 12'b0_000_01100110;
	12'b0_010_10000010 : r_w_inv <= 12'b0_000_01100110;
	12'b0_010_10000011 : r_w_inv <= 12'b0_000_01100110;
	12'b0_010_10000100 : r_w_inv <= 12'b0_000_01100110;
	12'b0_010_10000101 : r_w_inv <= 12'b0_000_01100110;
	12'b0_010_10000110 : r_w_inv <= 12'b0_000_01100101;
	12'b0_010_10000111 : r_w_inv <= 12'b0_000_01100101;
	12'b0_010_10001000 : r_w_inv <= 12'b0_000_01100101;
	12'b0_010_10001001 : r_w_inv <= 12'b0_000_01100101;
	12'b0_010_10001010 : r_w_inv <= 12'b0_000_01100101;
	12'b0_010_10001011 : r_w_inv <= 12'b0_000_01100101;
	12'b0_010_10001100 : r_w_inv <= 12'b0_000_01100101;
	12'b0_010_10001101 : r_w_inv <= 12'b0_000_01100100;
	12'b0_010_10001110 : r_w_inv <= 12'b0_000_01100100;
	12'b0_010_10001111 : r_w_inv <= 12'b0_000_01100100;
	12'b0_010_10010000 : r_w_inv <= 12'b0_000_01100100;
	12'b0_010_10010001 : r_w_inv <= 12'b0_000_01100100;
	12'b0_010_10010010 : r_w_inv <= 12'b0_000_01100100;
	12'b0_010_10010011 : r_w_inv <= 12'b0_000_01100011;
	12'b0_010_10010100 : r_w_inv <= 12'b0_000_01100011;
	12'b0_010_10010101 : r_w_inv <= 12'b0_000_01100011;
	12'b0_010_10010110 : r_w_inv <= 12'b0_000_01100011;
	12'b0_010_10010111 : r_w_inv <= 12'b0_000_01100011;
	12'b0_010_10011000 : r_w_inv <= 12'b0_000_01100011;
	12'b0_010_10011001 : r_w_inv <= 12'b0_000_01100011;
	12'b0_010_10011010 : r_w_inv <= 12'b0_000_01100010;
	12'b0_010_10011011 : r_w_inv <= 12'b0_000_01100010;
	12'b0_010_10011100 : r_w_inv <= 12'b0_000_01100010;
	12'b0_010_10011101 : r_w_inv <= 12'b0_000_01100010;
	12'b0_010_10011110 : r_w_inv <= 12'b0_000_01100010;
	12'b0_010_10011111 : r_w_inv <= 12'b0_000_01100010;
	12'b0_010_10100000 : r_w_inv <= 12'b0_000_01100010;
	12'b0_010_10100001 : r_w_inv <= 12'b0_000_01100001;
	12'b0_010_10100010 : r_w_inv <= 12'b0_000_01100001;
	12'b0_010_10100011 : r_w_inv <= 12'b0_000_01100001;
	12'b0_010_10100100 : r_w_inv <= 12'b0_000_01100001;
	12'b0_010_10100101 : r_w_inv <= 12'b0_000_01100001;
	12'b0_010_10100110 : r_w_inv <= 12'b0_000_01100001;
	12'b0_010_10100111 : r_w_inv <= 12'b0_000_01100001;
	12'b0_010_10101000 : r_w_inv <= 12'b0_000_01100000;
	12'b0_010_10101001 : r_w_inv <= 12'b0_000_01100000;
	12'b0_010_10101010 : r_w_inv <= 12'b0_000_01100000;
	12'b0_010_10101011 : r_w_inv <= 12'b0_000_01100000;
	12'b0_010_10101100 : r_w_inv <= 12'b0_000_01100000;
	12'b0_010_10101101 : r_w_inv <= 12'b0_000_01100000;
	12'b0_010_10101110 : r_w_inv <= 12'b0_000_01100000;
	12'b0_010_10101111 : r_w_inv <= 12'b0_000_01011111;
	12'b0_010_10110000 : r_w_inv <= 12'b0_000_01011111;
	12'b0_010_10110001 : r_w_inv <= 12'b0_000_01011111;
	12'b0_010_10110010 : r_w_inv <= 12'b0_000_01011111;
	12'b0_010_10110011 : r_w_inv <= 12'b0_000_01011111;
	12'b0_010_10110100 : r_w_inv <= 12'b0_000_01011111;
	12'b0_010_10110101 : r_w_inv <= 12'b0_000_01011111;
	12'b0_010_10110110 : r_w_inv <= 12'b0_000_01011110;
	12'b0_010_10110111 : r_w_inv <= 12'b0_000_01011110;
	12'b0_010_10111000 : r_w_inv <= 12'b0_000_01011110;
	12'b0_010_10111001 : r_w_inv <= 12'b0_000_01011110;
	12'b0_010_10111010 : r_w_inv <= 12'b0_000_01011110;
	12'b0_010_10111011 : r_w_inv <= 12'b0_000_01011110;
	12'b0_010_10111100 : r_w_inv <= 12'b0_000_01011110;
	12'b0_010_10111101 : r_w_inv <= 12'b0_000_01011101;
	12'b0_010_10111110 : r_w_inv <= 12'b0_000_01011101;
	12'b0_010_10111111 : r_w_inv <= 12'b0_000_01011101;
	12'b0_010_11000000 : r_w_inv <= 12'b0_000_01011101;
	12'b0_010_11000001 : r_w_inv <= 12'b0_000_01011101;
	12'b0_010_11000010 : r_w_inv <= 12'b0_000_01011101;
	12'b0_010_11000011 : r_w_inv <= 12'b0_000_01011101;
	12'b0_010_11000100 : r_w_inv <= 12'b0_000_01011101;
	12'b0_010_11000101 : r_w_inv <= 12'b0_000_01011100;
	12'b0_010_11000110 : r_w_inv <= 12'b0_000_01011100;
	12'b0_010_11000111 : r_w_inv <= 12'b0_000_01011100;
	12'b0_010_11001000 : r_w_inv <= 12'b0_000_01011100;
	12'b0_010_11001001 : r_w_inv <= 12'b0_000_01011100;
	12'b0_010_11001010 : r_w_inv <= 12'b0_000_01011100;
	12'b0_010_11001011 : r_w_inv <= 12'b0_000_01011100;
	12'b0_010_11001100 : r_w_inv <= 12'b0_000_01011100;
	12'b0_010_11001101 : r_w_inv <= 12'b0_000_01011011;
	12'b0_010_11001110 : r_w_inv <= 12'b0_000_01011011;
	12'b0_010_11001111 : r_w_inv <= 12'b0_000_01011011;
	12'b0_010_11010000 : r_w_inv <= 12'b0_000_01011011;
	12'b0_010_11010001 : r_w_inv <= 12'b0_000_01011011;
	12'b0_010_11010010 : r_w_inv <= 12'b0_000_01011011;
	12'b0_010_11010011 : r_w_inv <= 12'b0_000_01011011;
	12'b0_010_11010100 : r_w_inv <= 12'b0_000_01011011;
	12'b0_010_11010101 : r_w_inv <= 12'b0_000_01011010;
	12'b0_010_11010110 : r_w_inv <= 12'b0_000_01011010;
	12'b0_010_11010111 : r_w_inv <= 12'b0_000_01011010;
	12'b0_010_11011000 : r_w_inv <= 12'b0_000_01011010;
	12'b0_010_11011001 : r_w_inv <= 12'b0_000_01011010;
	12'b0_010_11011010 : r_w_inv <= 12'b0_000_01011010;
	12'b0_010_11011011 : r_w_inv <= 12'b0_000_01011010;
	12'b0_010_11011100 : r_w_inv <= 12'b0_000_01011010;
	12'b0_010_11011101 : r_w_inv <= 12'b0_000_01011001;
	12'b0_010_11011110 : r_w_inv <= 12'b0_000_01011001;
	12'b0_010_11011111 : r_w_inv <= 12'b0_000_01011001;
	12'b0_010_11100000 : r_w_inv <= 12'b0_000_01011001;
	12'b0_010_11100001 : r_w_inv <= 12'b0_000_01011001;
	12'b0_010_11100010 : r_w_inv <= 12'b0_000_01011001;
	12'b0_010_11100011 : r_w_inv <= 12'b0_000_01011001;
	12'b0_010_11100100 : r_w_inv <= 12'b0_000_01011001;
	12'b0_010_11100101 : r_w_inv <= 12'b0_000_01011000;
	12'b0_010_11100110 : r_w_inv <= 12'b0_000_01011000;
	12'b0_010_11100111 : r_w_inv <= 12'b0_000_01011000;
	12'b0_010_11101000 : r_w_inv <= 12'b0_000_01011000;
	12'b0_010_11101001 : r_w_inv <= 12'b0_000_01011000;
	12'b0_010_11101010 : r_w_inv <= 12'b0_000_01011000;
	12'b0_010_11101011 : r_w_inv <= 12'b0_000_01011000;
	12'b0_010_11101100 : r_w_inv <= 12'b0_000_01011000;
	12'b0_010_11101101 : r_w_inv <= 12'b0_000_01011000;
	12'b0_010_11101110 : r_w_inv <= 12'b0_000_01010111;
	12'b0_010_11101111 : r_w_inv <= 12'b0_000_01010111;
	12'b0_010_11110000 : r_w_inv <= 12'b0_000_01010111;
	12'b0_010_11110001 : r_w_inv <= 12'b0_000_01010111;
	12'b0_010_11110010 : r_w_inv <= 12'b0_000_01010111;
	12'b0_010_11110011 : r_w_inv <= 12'b0_000_01010111;
	12'b0_010_11110100 : r_w_inv <= 12'b0_000_01010111;
	12'b0_010_11110101 : r_w_inv <= 12'b0_000_01010111;
	12'b0_010_11110110 : r_w_inv <= 12'b0_000_01010110;
	12'b0_010_11110111 : r_w_inv <= 12'b0_000_01010110;
	12'b0_010_11111000 : r_w_inv <= 12'b0_000_01010110;
	12'b0_010_11111001 : r_w_inv <= 12'b0_000_01010110;
	12'b0_010_11111010 : r_w_inv <= 12'b0_000_01010110;
	12'b0_010_11111011 : r_w_inv <= 12'b0_000_01010110;
	12'b0_010_11111100 : r_w_inv <= 12'b0_000_01010110;
	12'b0_010_11111101 : r_w_inv <= 12'b0_000_01010110;
	12'b0_010_11111110 : r_w_inv <= 12'b0_000_01010110;
	12'b0_010_11111111 : r_w_inv <= 12'b0_000_01010101;
	12'b0_011_00000000 : r_w_inv <= 12'b0_000_01010101;
	12'b0_011_00000001 : r_w_inv <= 12'b0_000_01010101;
	12'b0_011_00000010 : r_w_inv <= 12'b0_000_01010101;
	12'b0_011_00000011 : r_w_inv <= 12'b0_000_01010101;
	12'b0_011_00000100 : r_w_inv <= 12'b0_000_01010101;
	12'b0_011_00000101 : r_w_inv <= 12'b0_000_01010101;
	12'b0_011_00000110 : r_w_inv <= 12'b0_000_01010101;
	12'b0_011_00000111 : r_w_inv <= 12'b0_000_01010101;
	12'b0_011_00001000 : r_w_inv <= 12'b0_000_01010100;
	12'b0_011_00001001 : r_w_inv <= 12'b0_000_01010100;
	12'b0_011_00001010 : r_w_inv <= 12'b0_000_01010100;
	12'b0_011_00001011 : r_w_inv <= 12'b0_000_01010100;
	12'b0_011_00001100 : r_w_inv <= 12'b0_000_01010100;
	12'b0_011_00001101 : r_w_inv <= 12'b0_000_01010100;
	12'b0_011_00001110 : r_w_inv <= 12'b0_000_01010100;
	12'b0_011_00001111 : r_w_inv <= 12'b0_000_01010100;
	12'b0_011_00010000 : r_w_inv <= 12'b0_000_01010100;
	12'b0_011_00010001 : r_w_inv <= 12'b0_000_01010011;
	12'b0_011_00010010 : r_w_inv <= 12'b0_000_01010011;
	12'b0_011_00010011 : r_w_inv <= 12'b0_000_01010011;
	12'b0_011_00010100 : r_w_inv <= 12'b0_000_01010011;
	12'b0_011_00010101 : r_w_inv <= 12'b0_000_01010011;
	12'b0_011_00010110 : r_w_inv <= 12'b0_000_01010011;
	12'b0_011_00010111 : r_w_inv <= 12'b0_000_01010011;
	12'b0_011_00011000 : r_w_inv <= 12'b0_000_01010011;
	12'b0_011_00011001 : r_w_inv <= 12'b0_000_01010011;
	12'b0_011_00011010 : r_w_inv <= 12'b0_000_01010011;
	12'b0_011_00011011 : r_w_inv <= 12'b0_000_01010010;
	12'b0_011_00011100 : r_w_inv <= 12'b0_000_01010010;
	12'b0_011_00011101 : r_w_inv <= 12'b0_000_01010010;
	12'b0_011_00011110 : r_w_inv <= 12'b0_000_01010010;
	12'b0_011_00011111 : r_w_inv <= 12'b0_000_01010010;
	12'b0_011_00100000 : r_w_inv <= 12'b0_000_01010010;
	12'b0_011_00100001 : r_w_inv <= 12'b0_000_01010010;
	12'b0_011_00100010 : r_w_inv <= 12'b0_000_01010010;
	12'b0_011_00100011 : r_w_inv <= 12'b0_000_01010010;
	12'b0_011_00100100 : r_w_inv <= 12'b0_000_01010010;
	12'b0_011_00100101 : r_w_inv <= 12'b0_000_01010001;
	12'b0_011_00100110 : r_w_inv <= 12'b0_000_01010001;
	12'b0_011_00100111 : r_w_inv <= 12'b0_000_01010001;
	12'b0_011_00101000 : r_w_inv <= 12'b0_000_01010001;
	12'b0_011_00101001 : r_w_inv <= 12'b0_000_01010001;
	12'b0_011_00101010 : r_w_inv <= 12'b0_000_01010001;
	12'b0_011_00101011 : r_w_inv <= 12'b0_000_01010001;
	12'b0_011_00101100 : r_w_inv <= 12'b0_000_01010001;
	12'b0_011_00101101 : r_w_inv <= 12'b0_000_01010001;
	12'b0_011_00101110 : r_w_inv <= 12'b0_000_01010001;
	12'b0_011_00101111 : r_w_inv <= 12'b0_000_01010000;
	12'b0_011_00110000 : r_w_inv <= 12'b0_000_01010000;
	12'b0_011_00110001 : r_w_inv <= 12'b0_000_01010000;
	12'b0_011_00110010 : r_w_inv <= 12'b0_000_01010000;
	12'b0_011_00110011 : r_w_inv <= 12'b0_000_01010000;
	12'b0_011_00110100 : r_w_inv <= 12'b0_000_01010000;
	12'b0_011_00110101 : r_w_inv <= 12'b0_000_01010000;
	12'b0_011_00110110 : r_w_inv <= 12'b0_000_01010000;
	12'b0_011_00110111 : r_w_inv <= 12'b0_000_01010000;
	12'b0_011_00111000 : r_w_inv <= 12'b0_000_01010000;
	12'b0_011_00111001 : r_w_inv <= 12'b0_000_01001111;
	12'b0_011_00111010 : r_w_inv <= 12'b0_000_01001111;
	12'b0_011_00111011 : r_w_inv <= 12'b0_000_01001111;
	12'b0_011_00111100 : r_w_inv <= 12'b0_000_01001111;
	12'b0_011_00111101 : r_w_inv <= 12'b0_000_01001111;
	12'b0_011_00111110 : r_w_inv <= 12'b0_000_01001111;
	12'b0_011_00111111 : r_w_inv <= 12'b0_000_01001111;
	12'b0_011_01000000 : r_w_inv <= 12'b0_000_01001111;
	12'b0_011_01000001 : r_w_inv <= 12'b0_000_01001111;
	12'b0_011_01000010 : r_w_inv <= 12'b0_000_01001111;
	12'b0_011_01000011 : r_w_inv <= 12'b0_000_01001111;
	12'b0_011_01000100 : r_w_inv <= 12'b0_000_01001110;
	12'b0_011_01000101 : r_w_inv <= 12'b0_000_01001110;
	12'b0_011_01000110 : r_w_inv <= 12'b0_000_01001110;
	12'b0_011_01000111 : r_w_inv <= 12'b0_000_01001110;
	12'b0_011_01001000 : r_w_inv <= 12'b0_000_01001110;
	12'b0_011_01001001 : r_w_inv <= 12'b0_000_01001110;
	12'b0_011_01001010 : r_w_inv <= 12'b0_000_01001110;
	12'b0_011_01001011 : r_w_inv <= 12'b0_000_01001110;
	12'b0_011_01001100 : r_w_inv <= 12'b0_000_01001110;
	12'b0_011_01001101 : r_w_inv <= 12'b0_000_01001110;
	12'b0_011_01001110 : r_w_inv <= 12'b0_000_01001101;
	12'b0_011_01001111 : r_w_inv <= 12'b0_000_01001101;
	12'b0_011_01010000 : r_w_inv <= 12'b0_000_01001101;
	12'b0_011_01010001 : r_w_inv <= 12'b0_000_01001101;
	12'b0_011_01010010 : r_w_inv <= 12'b0_000_01001101;
	12'b0_011_01010011 : r_w_inv <= 12'b0_000_01001101;
	12'b0_011_01010100 : r_w_inv <= 12'b0_000_01001101;
	12'b0_011_01010101 : r_w_inv <= 12'b0_000_01001101;
	12'b0_011_01010110 : r_w_inv <= 12'b0_000_01001101;
	12'b0_011_01010111 : r_w_inv <= 12'b0_000_01001101;
	12'b0_011_01011000 : r_w_inv <= 12'b0_000_01001101;
	12'b0_011_01011001 : r_w_inv <= 12'b0_000_01001100;
	12'b0_011_01011010 : r_w_inv <= 12'b0_000_01001100;
	12'b0_011_01011011 : r_w_inv <= 12'b0_000_01001100;
	12'b0_011_01011100 : r_w_inv <= 12'b0_000_01001100;
	12'b0_011_01011101 : r_w_inv <= 12'b0_000_01001100;
	12'b0_011_01011110 : r_w_inv <= 12'b0_000_01001100;
	12'b0_011_01011111 : r_w_inv <= 12'b0_000_01001100;
	12'b0_011_01100000 : r_w_inv <= 12'b0_000_01001100;
	12'b0_011_01100001 : r_w_inv <= 12'b0_000_01001100;
	12'b0_011_01100010 : r_w_inv <= 12'b0_000_01001100;
	12'b0_011_01100011 : r_w_inv <= 12'b0_000_01001100;
	12'b0_011_01100100 : r_w_inv <= 12'b0_000_01001100;
	12'b0_011_01100101 : r_w_inv <= 12'b0_000_01001011;
	12'b0_011_01100110 : r_w_inv <= 12'b0_000_01001011;
	12'b0_011_01100111 : r_w_inv <= 12'b0_000_01001011;
	12'b0_011_01101000 : r_w_inv <= 12'b0_000_01001011;
	12'b0_011_01101001 : r_w_inv <= 12'b0_000_01001011;
	12'b0_011_01101010 : r_w_inv <= 12'b0_000_01001011;
	12'b0_011_01101011 : r_w_inv <= 12'b0_000_01001011;
	12'b0_011_01101100 : r_w_inv <= 12'b0_000_01001011;
	12'b0_011_01101101 : r_w_inv <= 12'b0_000_01001011;
	12'b0_011_01101110 : r_w_inv <= 12'b0_000_01001011;
	12'b0_011_01101111 : r_w_inv <= 12'b0_000_01001011;
	12'b0_011_01110000 : r_w_inv <= 12'b0_000_01001010;
	12'b0_011_01110001 : r_w_inv <= 12'b0_000_01001010;
	12'b0_011_01110010 : r_w_inv <= 12'b0_000_01001010;
	12'b0_011_01110011 : r_w_inv <= 12'b0_000_01001010;
	12'b0_011_01110100 : r_w_inv <= 12'b0_000_01001010;
	12'b0_011_01110101 : r_w_inv <= 12'b0_000_01001010;
	12'b0_011_01110110 : r_w_inv <= 12'b0_000_01001010;
	12'b0_011_01110111 : r_w_inv <= 12'b0_000_01001010;
	12'b0_011_01111000 : r_w_inv <= 12'b0_000_01001010;
	12'b0_011_01111001 : r_w_inv <= 12'b0_000_01001010;
	12'b0_011_01111010 : r_w_inv <= 12'b0_000_01001010;
	12'b0_011_01111011 : r_w_inv <= 12'b0_000_01001010;
	12'b0_011_01111100 : r_w_inv <= 12'b0_000_01001001;
	12'b0_011_01111101 : r_w_inv <= 12'b0_000_01001001;
	12'b0_011_01111110 : r_w_inv <= 12'b0_000_01001001;
	12'b0_011_01111111 : r_w_inv <= 12'b0_000_01001001;
	12'b0_011_10000000 : r_w_inv <= 12'b0_000_01001001;
	12'b0_011_10000001 : r_w_inv <= 12'b0_000_01001001;
	12'b0_011_10000010 : r_w_inv <= 12'b0_000_01001001;
	12'b0_011_10000011 : r_w_inv <= 12'b0_000_01001001;
	12'b0_011_10000100 : r_w_inv <= 12'b0_000_01001001;
	12'b0_011_10000101 : r_w_inv <= 12'b0_000_01001001;
	12'b0_011_10000110 : r_w_inv <= 12'b0_000_01001001;
	12'b0_011_10000111 : r_w_inv <= 12'b0_000_01001001;
	12'b0_011_10001000 : r_w_inv <= 12'b0_000_01001001;
	12'b0_011_10001001 : r_w_inv <= 12'b0_000_01001000;
	12'b0_011_10001010 : r_w_inv <= 12'b0_000_01001000;
	12'b0_011_10001011 : r_w_inv <= 12'b0_000_01001000;
	12'b0_011_10001100 : r_w_inv <= 12'b0_000_01001000;
	12'b0_011_10001101 : r_w_inv <= 12'b0_000_01001000;
	12'b0_011_10001110 : r_w_inv <= 12'b0_000_01001000;
	12'b0_011_10001111 : r_w_inv <= 12'b0_000_01001000;
	12'b0_011_10010000 : r_w_inv <= 12'b0_000_01001000;
	12'b0_011_10010001 : r_w_inv <= 12'b0_000_01001000;
	12'b0_011_10010010 : r_w_inv <= 12'b0_000_01001000;
	12'b0_011_10010011 : r_w_inv <= 12'b0_000_01001000;
	12'b0_011_10010100 : r_w_inv <= 12'b0_000_01001000;
	12'b0_011_10010101 : r_w_inv <= 12'b0_000_01000111;
	12'b0_011_10010110 : r_w_inv <= 12'b0_000_01000111;
	12'b0_011_10010111 : r_w_inv <= 12'b0_000_01000111;
	12'b0_011_10011000 : r_w_inv <= 12'b0_000_01000111;
	12'b0_011_10011001 : r_w_inv <= 12'b0_000_01000111;
	12'b0_011_10011010 : r_w_inv <= 12'b0_000_01000111;
	12'b0_011_10011011 : r_w_inv <= 12'b0_000_01000111;
	12'b0_011_10011100 : r_w_inv <= 12'b0_000_01000111;
	12'b0_011_10011101 : r_w_inv <= 12'b0_000_01000111;
	12'b0_011_10011110 : r_w_inv <= 12'b0_000_01000111;
	12'b0_011_10011111 : r_w_inv <= 12'b0_000_01000111;
	12'b0_011_10100000 : r_w_inv <= 12'b0_000_01000111;
	12'b0_011_10100001 : r_w_inv <= 12'b0_000_01000111;
	12'b0_011_10100010 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10100011 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10100100 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10100101 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10100110 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10100111 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10101000 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10101001 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10101010 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10101011 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10101100 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10101101 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10101110 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10101111 : r_w_inv <= 12'b0_000_01000110;
	12'b0_011_10110000 : r_w_inv <= 12'b0_000_01000101;
	12'b0_011_10110001 : r_w_inv <= 12'b0_000_01000101;
	12'b0_011_10110010 : r_w_inv <= 12'b0_000_01000101;
	12'b0_011_10110011 : r_w_inv <= 12'b0_000_01000101;
	12'b0_011_10110100 : r_w_inv <= 12'b0_000_01000101;
	12'b0_011_10110101 : r_w_inv <= 12'b0_000_01000101;
	12'b0_011_10110110 : r_w_inv <= 12'b0_000_01000101;
	12'b0_011_10110111 : r_w_inv <= 12'b0_000_01000101;
	12'b0_011_10111000 : r_w_inv <= 12'b0_000_01000101;
	12'b0_011_10111001 : r_w_inv <= 12'b0_000_01000101;
	12'b0_011_10111010 : r_w_inv <= 12'b0_000_01000101;
	12'b0_011_10111011 : r_w_inv <= 12'b0_000_01000101;
	12'b0_011_10111100 : r_w_inv <= 12'b0_000_01000101;
	12'b0_011_10111101 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_10111110 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_10111111 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_11000000 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_11000001 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_11000010 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_11000011 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_11000100 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_11000101 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_11000110 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_11000111 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_11001000 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_11001001 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_11001010 : r_w_inv <= 12'b0_000_01000100;
	12'b0_011_11001011 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11001100 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11001101 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11001110 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11001111 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11010000 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11010001 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11010010 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11010011 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11010100 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11010101 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11010110 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11010111 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11011000 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11011001 : r_w_inv <= 12'b0_000_01000011;
	12'b0_011_11011010 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11011011 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11011100 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11011101 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11011110 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11011111 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11100000 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11100001 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11100010 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11100011 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11100100 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11100101 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11100110 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11100111 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11101000 : r_w_inv <= 12'b0_000_01000010;
	12'b0_011_11101001 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11101010 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11101011 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11101100 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11101101 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11101110 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11101111 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11110000 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11110001 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11110010 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11110011 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11110100 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11110101 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11110110 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11110111 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11111000 : r_w_inv <= 12'b0_000_01000001;
	12'b0_011_11111001 : r_w_inv <= 12'b0_000_01000000;
	12'b0_011_11111010 : r_w_inv <= 12'b0_000_01000000;
	12'b0_011_11111011 : r_w_inv <= 12'b0_000_01000000;
	12'b0_011_11111100 : r_w_inv <= 12'b0_000_01000000;
	12'b0_011_11111101 : r_w_inv <= 12'b0_000_01000000;
	12'b0_011_11111110 : r_w_inv <= 12'b0_000_01000000;
	12'b0_011_11111111 : r_w_inv <= 12'b0_000_01000000;
	12'b0_100_00000000 : r_w_inv <= 12'b0_000_01000000;
	default   : r_w_inv <= 12'd1;
 endcase;
end
endmodule